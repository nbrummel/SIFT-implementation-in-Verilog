XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}u�V%.֐P�7�G���؁w�w��?�d��|��ح;A�t��v���l$�8�h�Snyl�s����_>����`�֠8�x���ܜXV�0ӟ�3؍�E�̶����%��U��������#�̊nB����C+b�OAs�"��~@/�Jb,p>^��Z^�?
�b7O�jz���y�2�yR���[h��S�͘��nefu�u�_72�8/��u���`D����Xs�q����P���<��n��`�#���"K�8Ar�Rf�\�<���������A~sb�;�N1Э/��sW����%	8�vk=�~�?��f䶁��]m�ܪ̥j�e�l���a��D#ڃLh	�Q�o�m�^�Fh������x��3a� �%��u��N۳[��IE> 0��g�T����/CmC��	�U�8��k��>�g�����9<��65W��7�^��ble1�)����%���m�n{K9�gx�P����,��r���_Aw����Et�aӿ>���eM%�pZ�g���yY
�t�j�U[�4 TT�Ƨ=2qE���)w'�:Ҋ�W��$e*�F���1Ј�N5�1���LS��α���>�7@���0o���I{��ԑLvc����,jxf�k�t���Gb�[���p��B�t�%`��7y�@%8�.�>	X�{�[9�n��U�2>,�� >N�Q8�ʀ��S�{V��K��F�D���ǀ���( gᢏ꯹�-e�B��,>90;�r#L�n�XlxVHYEB    fa00    1ca0�����?�^u��+�JG��F�����x��I'P��(R�l���'x=�WH�����7��3v5u�Qf�1�������6�k� �C�0U;��e��T\���k+!�����7�u�����%Hm��O1�<k�t�ݙ�#���nK\e�v��k��X��V�H����m]Q�K�MJ�Y��B�֚M�(B	�m�!��R�c�jǕ�rűc6���UQ���������q��܀�TtB��aᶉR��S�BAU����O����Sp�8��t^ß�����D>D�o�J�>�j��rUj���J�o�ۖmX�Q���y��TG%Bp�>���Y?;ej\��X�:F3D=t�"�a:�f�M�����`��E����S�P��O��������\a�9b�D�Ӫ� ��� >O#{Y��yU�#ݳO��������P������!ħ���Ufk��1A*:�OIQ��YoH�@���0�1VhNՒ�ܫ���f��D( �\�d��8d��

��c�q�:�ۼq�$v��{X�oz<1������W)t((��<�ix���Z�hS�fQE�2�-���_�幎f"���F�e�y��R��y���+l ĎtA�ʗ��Kx��%�O�p裀 8�����Xq���.MOQ%���ٮ8W=Ҁ���i�DK�Z.����p�$����E��ٝ'g}��u����ʟ0E{!�T#w�/6�H��|I��]C��1Y��^�/d�]U'�3\B�p☽��Q�u�N�}'a]������uL���+�3��w͖�R�حX�N�;G�7H��5�3SFw��]�1�u��L���lQ�ᑌ��f_Lao����Ds��/��)�G�5F%��3i����Tr��X��k���F��/w��ɤޠ~��͓{��S.+�M+����,��3$���2|������O'3��E��'�%�Rr�0?���V��/���N���ԐPɃ��i߶l4��iۯ&;.�,{iM���mP�M:��F;�`���#���52�3@�-��2�M�y 6���]v�8��7��_�{��;f_]
W��l�Ju�t��*#^� U����Ē7�Yb{pll0g��ȍ�~��*�ҥ�I(]�{Rn�&ԋ��D]��'Fz��=�'��N�|w��#�T��s�������nyF1 XZ9��G(��.�j�M�߅��WI+ܐ�`��w�&̼pn�LM�ʽyD#�a8R�g�>.p�2��M�[�}��<��Y]N5�[����(��2`�C�m���T�O"�\������/[�ނ�0o-��5A�i/,�h��r���7|�;Ω�knq�[Ն�z-��y�d�U�;R)��L|(u^[����-$5�J���&�6����r��6I�m�ЭB��V˾? 8"�ЏҸu�) �-Jcʨ	pl�"_����w��\�N]#�'�����+��8Ϳ���֯��~tS�ųbB�?al����鷗ِw�1�������pQ!
�s	{% ��K`�tP:��\4rm���8.����0<X�ڈ嘇�g]��|��/o q�6��!�Y��c:��dorq���BvR��-������}t�T 38�V�4X%�f���N������W�ҵKxf�H���#���L�K! �x]��� L�W/k8�� �ek1)8,�,
b��5X����P]��sw���t�M�.�i�t<�wy����P/��J�[�������>���Y��,!x��\47���jN��b���ǵ�Z���#�c��1��C�-����7(<2�T�m�Xd]�[�{l�!k�=���m��F�l7l��W[m�.�ih���g���O�qP"�K��B�ؽ���X�uP!�W�j�`^O��y��[�j&98�u�>VG37�s�pq��e�"H�%�E���������Y}�YEMn����8�GQq�Ӳ�޶��>��s�bM�'�ֳU���Y��@?�`�����[i�0�9^�t����0.�{�$<���
i��\�"e8����6��kQ.�]g������.��×%��R�+�ѳaJ�i���]Ya����#ـ0(�S�zN�n.P(�ٖ�5�𛿘�'�}Vq^g=#�q�R���nM��T�ܗ�n�o[j
�� ����!(��
�(|��"�=P�}���K������<������Q	<��w��?���]�c����]�k�&��!H�j���훗T�}���"PU�7�#V�$����3z�pm�f+���v�?0��[Vn���C�m���b�f��L��Wr���a���X����z�ר���ko� `��U���i8��7r��h��Ac}��,�V1�T�5:�p/D�O(?�lU��'P�e�k�M�wO�Ô���E�~�+#�w�ܪ|⵾���z��������A��������#M����$t�j��4�G�!�@=2�� cɿU%�>Մ�&.�Mq+�7H^=&?�"� l~+'ﶘr�r�hO+�{-�=��v���=�7|��',~� T�e�Z9r�b)5�9�:/rB�[�}Rx�)#f+_�	)������gg�s*�TR2�3[w�~�a���1�~w�pg;�¥GIj���,��d��P>�U�gˬ�P� ������6���-���	iTO� ��k���fJ�������$�C���[eWm�T#���:���J�nɟ���_�*H�~�_k��*\�kPP}g�>)���ۮ��6��|��8jc�3�/:�bF,�N<"fc��2qv]:rg��H�������<�G��N@�C��][��N4σ_l��h�_A����$r����DE]�������ʆ�	3^���&�*�.yL"W��\d����?�<�D��,;�[��Ջ<���+ٸ��і�պP��������˽�cݵ���:î�(�@׼[Ph좯��踼�'P�W��jUy��4�[��'{o�qa��L�E8O�^�����p�� �[�G/y,�����]=�6��Y�W�Z�[vY���M3��e���jЄg����Ĺߝ�A�K<����j��n���f��g3�3�O\��P�j���ΨB��������(O㴊��Ӧ�E7�6u$K�@��Z{��ȍ�x ���{���-��u��!��L R�hwfA-�Dk�{�:s|��|��!Cwǃz�Q69���ϋmS��6��s�Ȅ�]X:A���!
U��K�p��5E2>a+iϼI�7�E��LMV�E�z�W��h�� ����n�n! F����OG��8S;T���k��M!�_T������p��g�7��&m@u�U[�t�����~a}�5maeT�1h}}�0h�=����U< ��HVݝ����7;��U�v*\��/��ٔR�]/�n�ڜq�{�jt:�ok��,�o��B�&� ��j�69%>��i�®ЃI�����[�)�x��������-�e�T���ć�a5#Ĺ`f�?�xp�oz�_/8�����t�	�Ď�- T"�H̀�7�ᯎ���r����Dv:%B�-���^h�d��_ ��͂4\f�Xv�`ym1k����=q���+��9�l�·2���C�>����7#b̶�4�d��y81�Y�a��ɲV��"x� �U����)�lѥ���C�k�2I<��H`�I�W�ڙt�92���/��|�Uш:������-����Q��Ӝd��U�-�����`{G=6K����+B���,�T�������@�[0�
6������5�L���zl7�� ټ�������Ĕu�fCv[I���ʹU�SR�D̍(�6o����;�^h��i C���Ddd6jb�DN�V�}����|Tq_n��F/&�����q�'�M̈��|���9����Q�����G��6������/�΃g��R����c���t�&�_�ZO�J
ooV+�*��hy��1ݥ�V�HE����(4��^Ɉ�Lg���[���c/��{�#�%�VP����������h�����q�{�k�h���K6���P�E��@d�|���^�轤�m@�Ȳd�U^B�Vs6�nO�^�!��-��0/��"�#�����_;	'B_���$����DG�|�hvY޹�ʕ�;I�UU��uq!^�eiϝ�_�#E�t-}���D.��<�K��$J�Q��P��,��N����zr���`�P0Y�+����TbkF�!��YDkQ+�)oV������!V�6���H4��`�GRH;��"��(Œ*VO��f���f����O�sY5f�ܘ��'b��H]X��̙�qSM�t�� �7Q,���Ʋ��Pv������#����A�n	oOr,�{h��	��=�!�|(�\}����A���� Eȵ�	*�a�p�"�}��{
?�+O<N�"�jU�V�z.�a�����R-���e��|p��)��h_&���g��Qf&_�t̐Կ�Q^+�$,A��)4�h�e �7�c�$O�~�����sYDG3;���YAh��<W(
��Â[���r���t�p.FZ=䢛�*�Y}�h����Ǜ��&�KC�����[5oSû�b�]7p�4�{��j��g��j��'��� ��9�%���c*w��MX�=@�w��iK����Ŭ���Y�q�^���B�p^I�-��4	��#u�Vݙ?��:��,w�0/���b�턺k&���$��
�?X��dJ6�&�0�aÎaM�t� zTSc�K����a�'�Z�7���xj����yC~P����[����ܣJ�?V����S���3�zި�Eߺ1��#��-:6�P%�vW�v~v�U��j���#j=�jq����%���R%��C/��7��;������tm��&î���[���1u�g�C�P��{��6���|˘ܭ��1�
U
s�f��j�����=SڡJik��P�4*��hs܌!l�;R��%��� �h���29[<��;v�i�+�]r��F�_;�%k�PC��,:��#�K�{`S��'WӟT��ʷ���&����TŞ���[П��ҷg>)5{�vfFe�W'un��ڭ��F.t�	D�#G	�AA�*M�(��X��,�ъ`:�5(�X�c�ٜnb�ܼ�C�4�?�Ќ�%ؐI��z�,��	#��Z�;^�ғ��j 4�^�;��0Y�i�?7�tc��:ZG\Z$w��m�=#��R�E�w�;�9���Ü���'X _�|PPͶ �H!e\ ���?���}8Τ�Kb���]	����{$Dݴmg�if��!A��z�b	�>^k�T)o\��_�$�)�����G6�%�by�p��?>ۏ�x�M�9q���9`�&:YF�;䌙Ď~�Gꛙ��$#`PJ5�3(����>��E8.J[�~Ԟ�"��^��5��-����N*AN����.�~)���1�0�G�4B2�!�����M�p,'���B�;=�r�d�(���_��ï�.�c���x���v���>�b���?Rh���8�5�U2�0'�sh����58�{/0U�~;vv@�RH�a1���",Bn�x3��r}j{�x�m��/*0��!X�7��=�Q���[?�uR�0��SI?"�F���&�Zz�E���Ί�n�/�U6tO��8�C<J|�я�!��_2��~!G�J�C��y���L]G4d?����3hs}�ڗ'F�+���ӑ�/��p*g���)�Ӣ�a>�>"l��}��BY�7	�d�K����FZ#�Q��*�=a��VT��y��m �%rOe��Q�m�ɉk4dR�zEly��Z63��/�/�z�]��p����d�r��7ݽކ�hE�b�rC�������&5 ~H1��e6
l8�)O�u�f��=��^~��t�r�rKv�c�Hqgj��8���U�9�F��%�2�	H��rDG��A%d�~�Fĺ�e�՘O���3�
�=��@b���0�p�Y���ӏ��"`��MD����t�4ώ�#��#�hrJb�tSP����d`���I~�h��gYn���oe�]CDf*����o�|�[����N��Zg	��hE!1Ɇ���_Iٿ�{���jfQ����#�J'��%g�zsi����m|3�Kv~C,�Y�E��P��L1�4����Z�o"MU
��{�2OX���	�v�(/��4O���#6������q�o DL'�a���`���۵��0PTi�[˽��
c�O�A�	�0O�&N�ff0���������k5��2hAJS����c�bg�J8������6�6����,�U�Q7	�xQ�(t�%u0���J�\GF�@�
��ƒ�Gm�{8����k�Ɯ1��nqS�c7; L0y [Y�v���o�Q���oE�u���K#,|~N5�s�|�!��%ɠ�;۸�\��%��݁�$�5h��W�m���ɎS��*4w��Z<�}ȧ`z8���U2�g9���Aqo���T��w���@����"��K
���CBQmi�~��۴��v8���)��A�mb����h�1`���ᜡi��ni��m+��~�]�h�H7峞Y1���}�W>�U'#���2}�u"-x*��54��6�č葝N;��5'n:����)dQ��2��>�uj��%ǌ���'ŗ��^��>���m��Q���,dhFqA�9*�1|h��\<)�n�|���el߾��Cn��a}>�l�91r�@B�E��芰�W	tq?�D�Ƽj�[�o�`.�)'��Ԏ?Mb�\����VC�!�|
�H������϶i�F���H�2:D:��n_}�\gCΆʽ�S�9sJ�7o���"�넃�����jٜG�\�	����ݸX����2�x���3L�WG������m��Ơ�xS���N�%�X�ӭ�DG[9r��pn�_��d8���W�z��A�"��"rd��Hr� ���˕�É@<7�����]��?���^�Q��~�\�Q߱�T"Du,f��5�e��,M"��kW*���O>^r�W�>����ȅ9zýb�}}<j��>�}�_ޮ%�;��!u�/[��tcE��ؤJ;��㙽��r�V� ���!��a�5�|�K�-��0�W�_�_��߻�hR��W�U�K(f�;���q�8�۶�XlxVHYEB    fa00     cf0YC�yz>�p�-�?TLt,��r^Y�<�4��F�Zt��a�ae�fإ�,��`�+���g�TYobSM�t���I
e��?�x���,�m �'�_-�gΡ.���5O�R�%�
���I.���{2�fB3����: g(�OK�� ~n0 �f��>�S�zy��I6�X�%�o�X�`,�]0�g� &�I�`e�� aS��4!qV�Eү�����z����~b��Oc��f�O��ߞ:��-rdq2�S֙T%{5���tq���*2�����ŏC�Y'O,唍��32�����qB��R�6,�S�U�zx�`w���&9�q����P�ȉ�1uϢHU4�H�#9�.bC;�)Ǳ���)�L�t'LL�T���m_S�Uف��E�}�T����w�KdJ�O�kó�&ٳ��6I�ך-6r��;��������+��踏���|d����ڶ����j�`'��Nb��i��ʏm=l��up����������L��#�r/v]{_�k�w��uzN�7�y[���#;<�*U�ju.��w��
s��w��u���,��Q�R �,��i����eb?H0�x�H|�,�U����^����?};���1V�7�hW+�zi)�}����k�=O^��1D��~ ���֝���!�`�4`I�2ݹ&��B}K�:�V���(OLꨗ��΍`�ݙ+hRP%{�Q���Wx�3�����?���&�|��~�Z33��;]�l�sl`�cN.|7j!&9��7J�����#��Ed��|U��к�L�8�pi6��y0X��\�R���jh����z������5�JE�pN�f��k���4{�H��N����U'̔�q�[v�"� �2�C�Ns�3c`�$F/i�N�[�MQ�F�#�P�pz���O�<��#�u	��>�J|go�!�4�m��
q��Ux|�3oO�b'j����^
��QUa��MBj�-��<r���<d�R�9S�Ia���<��$�NC�ZM�M=�#��=E��k���`���VO|5��!�n�B?�f�ΌҴ�gP%�b2�r՛����O�9��9�����@]�_�/r����&f��D�O{"MT9k}ז�v�rR�
����,�S�6�F����ҩ��	csI,O�3%�{;�
��pgڙ̃��6��)�"�E�\��E?�����hƾ;@���<sZ)��h�	Y4��m��z�0Z�����mLy�r6BZɢ��/�j�,�����wc��{+UgwQX��͝�* i?z��S���,hm�g��:֋Cޚ����V�%4����.)����N��N�$�g���zFd9~^�7��9�E-� u�@)����Uv�f�o��c.3.���%�-�C�D/	f&ݹ�3q��I����ﻹ�+��Zv��(�͚q,A�>�����P)�����|��%e2�K�F�u����>�GP��1�/�S_�+D�7�x�#�G�5D#L:�%���gɣ�����L��V�@���ͱ��_�:�57�ޮv�S�X(""�|��$�8b�B9���>�A��^+�n�,�p���a�;�i��c2�.������<��Bt�%#�-��ҙ�(�� ���UXS�$��zq�E�� �5ވ��MD�,���6���h�)4?��`J�?���|��%�V=���)���E��Ksv��2��FT���90J����,jd08���1�,�X
Ժ�q���J�J��4��%�d��_u��X��*�9�e;r�H��U?��Y��uj�5��Wm?}���m}��!Ɖ�̣�:��K��,Y�dgbkV�<�Qz���]Z�X+6<��^���n�v6{d[�P �.�>6QS�BB���d����kE���-�2}4�7
�)�$6���=N�>j1�'����g��� 1�f�s;8_�x��X��Z��p+�5g�Jɗ��;B4)H�vT��܂�7N�]�VD���aH>��?�[�Zá�dY�r#R y��z�X<�}Q����uż���D�IT�U1��ĳw�Y�DnCf�a7ֲ����!�9w׫	���kyF+�ʢ�@4坲Kg�ĩk5��){3�}v7Rx����n�*a�gÅ��K����m�>�XR�����d+@|gV��+�;�Ȧ��Z�P��de^�ܒ��B�f�#ԧ5��dQ7��ۍv��>t��ƁHk��|F'~�iHM��3��Knd�e?�FB� �Ow�ā�$<���k��LE1_���XI�w���0�vϰ	���y��3Ljg&Ր��N
�$��%U\�(q���;�=�ט�,��$�C��;�R��E�u
�d���y{uO��g�|P���kt�m}|R��Cqj�4��y�[�R���/�ZA�imj��K���j�>�veID�Ϸ��eFJ����@G?��r\\4��j�C1��*����,�2�'� �M����a�l݊A�f�[-!$"���]����,�ζB��Hłiߘ�����6�,���m^}V(,���,GM���]�
v`E̩�� 5�RW�n*[Ze���aE�����[�իO�G��i&�9�z`1?L��:�����5��t��^l��WJ�^�y.E�z���@��@�m\{pH>P ��{�o�֔�j
���bW����v�C$��=�T���,gư�s����L��t���B�.�T��z�D�7�<��y|�ۊ>A�w?�TۯU��J`�w�끶i%�n�VU�\�TRU:��;0�����Ic�e/�X>,<pf�d���G��S&x�xg�7� G�>ߪei&��8f8�\��湃`���Z	喂�^�?�x�w#�����U�dG����p�\;\��
�ɞ��
��5�_i��#�l哃��b:�K�hj���N@����0NfB��r>Ƴ��5�cf���,\��Xz\'��v��N�����C	kSƖ�6 ��w�@]wޚ6�U�r��`��/�rR�c�%N�����!5�Z�?��"v��pO+Z��W%�.z�7�d�Y�'Trb��Z��;�����FZs\\ݻ�4����9,X�}��B�3;Z��F��Uz��Ȥ�Rz��?QlHI�\B#��v6��5o�>�Y������V�갣P6i]z�h`ɦy#v� o��m��R���(d�X���-"��nm!��
�z��j$��:ļ��,��6ߤ�� ԔY�&��se=�9E�Э�S<�uI�S��l�B!�r��3�
[��XlxVHYEB    3981     4d0���Zz��e�sC���HS� �3�;Ψ�mB�ē����{��-Y�񀐻|�@y�I ݷŬ�����2�8�8�ѥ��p��;�����P8�&�5����|�h%��G�,�v�ܪoڕ2LM�u�\ D6j�X7!���H��6��KV\5�yS��M�ģ9w�ڡu5��Ij�\��R'�㮞Ȥ|���g"r �������JV��N�	�ia�^��P��ˍD�E�.����K��@�a���K�\��m�f�G�Z��U������^uXӭf<N�3�q�!�b��R4@/�'�K_NY`H��BS��B���kF��i>�P���>���f�'{�#��0���r�`{�_��I��̖��ۮc�*��1ё��)[2���h���	��	y��!��3�kZ�X ���ZJ�{k�j���(N\Ե��	g��!���|�vh�o�H�q;v��"իv	|� ���x}ȶr���9o��ǻ8?Z{H)��֚$R�{�>������Ѣ�zI��0�q )��Fh��U��	��u�=��Q�����d�!	���t/�J�r\��L��gI����D#F�y����MU��G�\X)<h�4��;t4���9(�%�a���=]q��	�L�ԸrS�FJh�G�Wyߒ��c
���&�����J����ck{w;��a�߹H�i�X&Y2�]�x��3C�ϭ����DIV{%�0�Kl����䮃�,|U��`�������_tQ_� �x*8|��8���|Hh�3s��?gh3��T��q�@Bz�2���ph�n��1]/�>?z�,Db���L4�f�̍�j�x��U�٩k�L���(F��f�xKy���7.�B���*F�/7�ur��'��+�����f�j�{�y��L�0x��C1��g�U��6)���J �#�e�7זho����{>�G!!V����kP|���9�4�ޫsR���3�~�`|Pf䔫� TN-2e=B+���PP{��.�����H�EVPk$�~�b!(T%���KU;���4u��t�jR0Uy�ѹ��	����Kȿ�~�L���v����bu��h:ă^eWcژ�P�S��O+ UEk\�⫬���:��Yg��B��yQq
�(�m����4���A��BU��-~(��Ӻ4p�m�s�oL�e�u�A��S�nJ�[5�K��S3�8bA���i]Q��&J