XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#W��	2�i=*�NU	P����~��K_���<��* jƭ���1;���Y?��R�Y��#RDo�BE`0�9M=轖��0sw���n(��g2%<�׮I��ZYϜ���к��Z������I�B��Ɛ<.dH�H1���y�B��*�D����pr�o�:�Pn�w�7�U�bn>���q�g�+��R��9h���F�6�0�� ����TH��A�;"ʕ�lt���Y�1~V���釀�H��\�}����c6�Ϛ����U����u���7&j^�Zh��[.閄�{���a�~/�a�|`�r*�>�u�\���/e��%�A	d��ūxf��h��#�|ԋ�,מ�>~�?&@��u	�Ս�:�3C��>��D�p; ����7T	ʀe_�7%|���7�qc��/(��ְ�w��u��=��b驩読/�uF�����7,��N���0�o��$��ʓ�Y�r�:���h�mG�������6@0��#���m��3��<�m]��3.u2�مl�4g�$�)Q�� �h��GA�d��C��7�e��Ǎ�A,D�����ED�,�
)F0��)�G\H�RdBe�fxC3�" 9ޣw���^���͖RA����?��1�R��Z����ޅ����ʺ5��v��2���"`^�q^��2r�J��p�(�ƻ*)�ʣ�e�����V5}4�>�?\�zt�����d��o��nhŁƱ̃�_��͵"F_7�P��,��$3C�D{���T׏/�i�XlxVHYEB    fa00    24c0�#��#���'���W�ڕ�QS��!|`r}��w�W���[2����:+FŖ$33m=4垗X�o����2yf	E��>^����Y�速PY
�#������^PW�z�;FOE�H�e�=��!���>KW�J�ҽ7�|j�#�HX�YP�w��'�[ɿZ�q������&LMj���/�4b��K�8��c�4��: ��e��jC�{�0Ta��p�h���l���ulH`]*��;!X�ԟ֜?r/B�\�<Fz׶�;�q�;읱���"���1�����8lAh��C��Eɝ��H xq�������a߱e)���ڌ�������2��+���oE�	F�f�e��Y&i�X�N�X~��t� �;�hܪB)6촅�Y^�^����$��ɧY�s��=�N���,��Y�ˍ�O��A���n ��[���
�	�~P��������c^M��!��)#ZDNH�%\�?����$g(5�P���,,Ƿ;Ptl����Y{}>���s�O3�5�o����`�""B��?(����\�|@���[ģ�{���5������sN-�b�x8r�����a0��\�����g˂1� CAcc)KD]������»x�R���&�Q��'�B���zL��Ux�Ϡ��w��2`xѳ�a�/�S���\a�}^��W��S],��������. n����5��3�S�SN
�j��<�:���j�"9@:_����Y��ΑM�����@�X�>DI_�y)o��~�9�Q#,���O]�2���>|�������-�Σ!����G�tnP�=�ʋ�$Ȫ\�0;��`ɜ"�����ه�Ah�]:�v+���߃�IҒ�b�2�;�����2�62�oYk��0�׹�\���	��/��o��zA7!�&��'�$�X!R�u�@G�S�a������
Vejgi���7>�>"������]�n'�E'��ji�
���
E�/��!��m	ңR����C�W���0����5ܴ��-F�63X4��_j�Ši���WP�ߟ�M��-A�!�5�4�ǁ��p�u���]�0?�px��� V?eu�j��k� �w뤧E��ɤ"l�7bh��0�E".����1�Oݽ�H�JGva��Xg4��NKrԮQ)���z1��ֲ.b�q�В�,���W�(niC�|�;�`�.¨s�V �Ӎ�e,�g��4�T!�%�(\�K"	ֻ?����eػ�P�c�����L����	��V]�W�Y�M�$(���;Q���m(]o���5#}��X	�ۇD���r�t�u�w�|�7���X;D�g{�]u4'\<���ԝ9/ksM�E \�1u���:ΏB���/=�@�d︺�ԣ;�n�	��q˙�/������[�a���������|� �9�{�&t!��c?�	�OW��=&�&|Ka��P�}���[1{����q��ߗ 3o*(�1z����<����m>�0�7ԎQ��.>�*�{W���1*���ჃqOHy�x�o?�λ ,���6��<�P��3v�����Y3-ڽeK�OA�y`3� �,��������b��ʞ��T�(ߣZ"d2h�5:�;��"&�k�Lz_��N�fS��S�Jd�� �Q�W��U�?��_��U}�ΖΣL}z�\�ll4s8S���\�}�,��`'j~��m�F���V�=:�_*rrhA�0lD�ա�ΐ�1Icۄ���7"�7$�Ib3.���
y7]hV�a���Y�vgИ���90��$��Q>ܽ�1�n�z���S�x�y�bN��I�ȫ8���#�&^�#��#dƗ�O��M��6���a��bF�q�b(f����WE
�R('@\��Sn�U�(]�MK�$�j<�*��	�z�v�������Ț��צ��"`��S���y"ͥ?4��%�mˋS�<���Gjþw���u�OID*�n�|��҃�h�,��T�7�D�8�f������o�Օ0o\�5�
�πv����N���>����9$13��j��;����SW�H�_����*�^*0^L���N9���E�]�YF%��C?z��XyĿSm;��ci2Z����nf���51D�����E6�"hK�>V<��%hZ���D�an
$`u}�߬i��PU�vpf�.�� ��Gk�j�A�����9��o4�9�Bosg�Ky��!Ɔ�jh
����6��1h>�$�5�Qg�b+���vD�Ħ�F����jǘvQ�=~+�1�U}K��X/z�h�����������1�9�>m�I��Z<�):֠U{�.�����/
����7��&����nor�In�/+�2�q%��b�q����?���.dR����1��aN��*�טּ85�	�������˘�+�$\1'��I��l�����n��dQ {�m}}���B�ӈ8�>2^eq,��j��л�	 �E0r�r�h�&�����h�����9���L((�u��;�U���k�w.l��U����ț�:�ET�X8�y��u_*"�\�L ��)s�N���m_pp�"�� 4�`����.�~^*�ɱ��g��W8\���y���)E̯������ͭ\��{; ��Ǣ�nG�g���b�Ϣ���,�?��_����!����Z*a}���8����e��W&<��ȉ���X@e2���x� >�Ɩ�V�֗��v_m�E/��i�(�䄐�$�7}J� ��r�����ɽpy�jF�0�Z�r9�,��� S��w"��+[i���()�*x2��:J�����d�`�;%��#��3��#����uY�G諪g��� ����#����[�"mnh"��Y�w\�����:�f�x"���w$��K�t5oe��s�%���� �Δ���X��ޞ�8d!n���z=�v[�:�5���x�Z]9��N� �=O���:�$ޟ��� �)�-N�~}�q#W���P$��1��_��/}�~B�9\p��8?��m���²��Ȧh�I��~X�рNV!����d[�-_n|��#���S�w���*!6'���������������DQ�:#s}:T�y��bUݾi��uM�6L�({��H3l[׬$(g�OY��ƚ�neC����އt��Ҡf�d��{�;z,���W����S!��9�������pǍ �s ������;!=b&�������n�ǔ���+����Q���ؿnO��V�ye�;燅=i��P�����Mk� (��|��j��*n�@���|0#b�ңO�d���*bU ������^�"�ʺ�1�����B�ʙ�`M�k j�L��>�m�!U����H�Bd���m���LV�ß��^4G���&�$��̠@����	�d�v�j��#>J�u$��u�� ����������T�Ӥ1�����S�/[�k	d�1h���T{�ƵfW���������ҳ���˧-�D�E~�ݝVt&�:w��wԖ�4�kAl�lJ��"�ל���d�M�:����]��۽� ����S]�B��[�E�XN�������#o:��6e�Cd�;�&��;��Ȕ��5z��c����� �qN�F�)Oi6b�F��㛪��x�Py}�`�#����9���J����D'�܄����f���x��cu����
lo�� ����d�PE�o�Ñ�Xm��cթ/��xf�C$g����4$�=,8a)!�
WA{�l ��AQ�G�����^���/���>���!X����}�I�*��cg-~�2kO6�w�6�%�<��jb!��Kn̢B��r�����a��!@�ڭ��EXH�Nb�u� >�ꅲi�)����n�m�"Y��H�S4��}��a����4� h���ެIw����M ���cE�2�*6,aU������Ԇ�x�qW|��_騑�o��Y�4�)�lp���5G� s�&G�U-���������7X��&pjLZ��`� ���:�9��\l�_�3`�5�6:Tc�8��*6�u�����R�z��z�a$���}��p��:IT{94�w
�6�r��:5���.>��̖s:���V�������>~hjir݇&9\�;|��b�z�"�ew�ݹ� �2h�Ub�Uc���,K����]C�5t������>1W�ý0�)_Ќl����(/��U'@0�����O�|�q>�i9|�4���:�m+޳4ǔC�*�TT���~�-��:���/iAk�J2s����Qū��>�D��n��!3�s��|�����G�x�3��C(09	����Z�W0~WM��YR`;���i�5^�@G�5�VM�p�c1
v�eA�P0��ґU�j�dkyF�?�
n�i�vA�'��}�K�a�~��v�qe�����U0�]���K��O�a&uo�U��˗4��a��	�6y<��λ�ā���$�$�+�Y����y���M��D������fE�c���G��(�sW�'P�m�����$�����;@��N�D�j?xL.�-^�� 6�����t2��l�ʛn���$9����N�hF9_s�)��^�Z%��c曾����NP��y��Z�z ���B ��8n�b�ާ���"�b�%]�lx̃�pCtg=gW�\S{�����7��޷�o�s�;���v�Ѵ�`懊MM�E�mМS��!���_Y<%Lk7��a�n��8�!��-����X�`�6Uᑠk|C�0,b�������>>�̖���߃�ǃj�}���6A?�]�`�3�C��-���~�n��Cs7�YP�f���y�r��GXhXʏCʹ?�[��WE��ē��d�=Z\��tiZ��Dݡ�[�v{K�� xb���7���[���Fg��U�M��*��٨�v�Qt�Ў��O�>An�>�z� �.��q��K�%��Օ��:&0�����T$@Lx��y�Y�`��I��(.���jp���*������2��sVl!��l n����,X�7��3�:A�B`��@9UÎj�`i]��#���"./`��if��<̗��xP��>%���P\���0
������	��k;S����xq�D}]+�r�Nmym�3�@^<k��u�%�L	P�d�xI��O@��M�ĉ�z�B�n�74���Pg7��a�G��T�߹I��5���䏨�mi|aY-·V���+7��ݨ�`�����}�w�Oʍ�rt��&Og�A�k�H~q�~CG����LH�-�t�k��vD�+��.�����{���$���R(�EV[�=�z$lY�����G���Az_�k�`2��y��Y��n�Ѽ��̔�>�u?z<녟�m!��΁�M�C����Coٱ��]�w��x�S��I�ɧ����oѸ�Li��&�X^'h>g#xX�x��9�]�"����r�/&�+q4�\�/h�D�_�԰qz-��r�,�U�w�5Ř�r����Z�Jky�8���>��޲f��fs����83��n9S~j��Bn D�Hǿ�״��{��~+n��M��P�����  Z\oL�w)�����~~�vV�e˪:�r| 
Իkr�t¹��M�ŁZ�'��Xp�$��Jv��M��yZ�?�4�DdЭ�ht٥B�;��.0R�u��)o�?oNC�)7Ȧ�?J��M:%�] �H,R|4V�M����V�Z|'��	�����)U���1�����9���
h����s� j�i�����.D[A��'��R��D���u���:P���N���X)���vVr�3!($���O6%�n'Rn}7pS�/	T-s��g�Wi���M$���2���$i@��6���8�X4~�+�����iv�\`N�*tК�t��<^D�ܘRI�On0�u�4���3��!]�eŴoIU��_>4���<���*cs�y��k�o�à[�Q�ra�*3��X���f����/�Kl�`��$,�[t}/wI0u��*^x�TL��`8N^����!�̪��9��� 3�<d�ɒ��,�^U,�=�ѯL�[�_�9P�u�B�x�7=�#g��Q�� m�|O9�vUw�>85��ȄF��l(�M;�.�	:�?�Q9n�[�ԅ���aIT��3&��W�<�@�w���s�d��-Up#��+���t�T�H0�p�M"H&�!z#��&�_<�?�fM4Y�Q�	݄Ƭ��?��bNP�0Ë�y�P��h�G��dh�[	�P���N]��%JOb�"�P{i��x���ؼ_���	����w+c郌�"��]�V�9�e-јN�H3�_�<�}S��M�Þ�J)JҺ�cc��I��}��=;3?�~��.p���L�R`f.����{`6i���ej 8On���s\ۙ�b�Ԃs�M�� JuSla�m��K���fQ�6ʭB�0�������p���8��j۸o���W�璲�>Y�g#o	�&u-&[{�U�����Q`����qO�(�ƫ�m�Ņ4�*Q"�EPMt�t�M-���M�����BǱ/uq��ֺ��O�$��D�A)a����$^��\��>\�8���0-��8�?цe�H��s��y l<b �����f(�f'R���u~-���`#q���i`+17�Z�C���3�>iɀ��Eǉ�ג��Q�&N�d>n�����Z�UB��(�jy��A� ����~')�J{\Z|Z���(�N��6	����^7+l�Q��y� ��x��x��g���6@��`h8lu�6�bY�A!���^0�M:*���:�Tڏd��oK�^����
�ݸ�[���S�6���4��M5B�/�	��0fI��itl� �/��r��%���X&ao�H�����R�
L�9|F�#�`!�#2���s�ƅ�3=�ߏ��DYd�{��� �X<�h�MH�;1���y��:��h�F���*4Ue����9>Ć��c2�+sW&��5���/�l����:��Sg�����bct.I��E�{�0F���O�v�x�P��@N�J���xN=���/�R�e���a�F�v���\�tG�]#E�_���b�9&���0�|�Fv�KWF��lm�#]���{n]�'/q̛�å�Q�a�@x
a�8���B@����,+����L
�pl���W��ȕ���k6��������r8W�8ݽg��yћ�X���{_5��q�S�)Յ��з��vO�������'O�*fv���&E@�-�#/�?@v�<M�[!G�|C��q�����]!2.���wJ��� t|ߞ$ ǤT��P��j��f�42�SU�3s6���]�H�z��}G��`#��i��.�5ǿ]�}E�����[�E�qD{�/�e��Eӭ�f�9�6B>�x�b�
D���,�}��Ŏ��؊8^0x��E�L����"�\Y�&�hZ�
�e�3ַMY�F��{e��
t�$:���Q°ǳ���g�<�,�]ĚݛoD�1���|&�
;| �7tq"��Ru�Y6my嫌�������畤��t�ݒ�̒%�*�$"�n�CQ1Mzx�Y#:�A~B	���if�\l�(���x!���p� ~`�\��4����3�[��]7��O���n�F�"kZ`ju��n�b;*�I����R�G���l���b`�f�6{\��_�Uh)�T*)��������	��V��S9=��O-��֍��r����L'>�9j[��:K+�8��k���;Έ���zp��$ǫq�95"���f�Q����0�Ԫn��ҋεx�cu�����ֆ�گ�*nȐ��� X�����:ކ��,i^ns���[�=uS��,U�#��lſ�����l�e�!T.��r���%��@���F%��!Wf�V9���x�gy��!2���D�-;G��O�x��E�5�N��V���uP�^Y�������u�����uAx�I�Zw��6���e�\c��u��X� ��R��N���9�y�������� ��7B{1Y3�`�d���g�FT����Ϗg�K�By8I�PؠB���H@}��ڤ١+`�I�/If_"�}_�`0�
�VC>9�z����9r��d£�l�?|�1D��S���M������-��i�>e��Ġ�R�*�_+���M�w8��5,0b�����=���{�^3�F�m`�x�X�к�8K,3��V^:AU�J,"!��K��%P������ҩ��B����]��jo���0��Ӧ�:>������BD�Úa�G3풀S<��~��'��dЏ����ݞ��?r/R/;̛�Qjriwq[>���7���B�r�S鵇����L�`��ؙ��qm{Y��]��y`�
� c�u��.�I4L��QRj=e	�R0�N���)tu�ͳ���ɡ���aO��/s7���*G0��C�|2T*h���ZmS�������:���C~}���0T����`��N2� O����,�$��u�o���E�W8��`��+ �U-��҈��Kԣl�4?a��������cm�$\�]��]o�VF�Z���a��j���'�I�����r��`�%��5ށbc�\�B��*)@�=�
*���G%���ּ�b�4�"	�p	��9u����_��A�1�gv�NB�t���y�u��bD�$8
�ocX�M��Gm��pq0Si�U.u櫴�N���O����G1�RV㤼�ϧ���t�*L�d�Ck?�]e8L9	��h	���%@�x=B��W��8:C�ѱ���&*Zú�AsN+�x��m�'"�$��+(�_��ٛ�~z�׍��Y�ܧ[��bmȀ���������R��>�n��[����J���Xbe������W=��VܱP�/ġǕ����6�X?�;!/4F�l�_U����>S+ԥ=�5����y�%�hɨ��0��2�U!�#��>t�D��K��b���i�
;}�����f�@0����q[;��x���c����]��(�� �S1߁�
�Oma
�\>��1����n~��Smrb�f8�=�X�����JXkK��)�	0#�N����@2�ã�l�H� 8�uw�j%I��?z� �e�U��#�tU��%��Xl������_,5`=��9������?*q�����53 ���u�bnpFM�i�נ�#�Iؤ���KG�~W],8��P�,�(73�����N�/��#�A�/��݌$��#������ߗf�P+�l0�M<Uq\��A0�c������d��-l�[U�񗺯�M��.XlxVHYEB    fa00    1e20Q�����֮�U�r�E�}g���wѲ�O��q�u!9�l�uH���� 6c���=���Q5q��ѹ�ų<H���󜪼��,ZXЍTR��x!�8�8A2�,�TJO��;��s2v��I\��hB���+|�@c��N��D��@�D���B��\:����&9�k��~b���\��j+x3Q�j���՘�d��;61/h��\(&�������Q��rR�U��CYE���3��B(�?��c�t�"fO�X�y:x�� ^�a�-�c/W��g	�\�M��ř�\�v�Q����k+KVh	���Kq^���V�,�9�t�uȋ��hȖ�d�<�-�������q��kyДhc��Ci}8֨w.�9��s���~x;�(a���]��I7-*�J�T�� ��I��/��}�0�.v��q��̤Q_��5��B��K%����Nfc L��!��N�	�-�.���s,����������ް���A��jw�������X{�Ȯli�g�|Qh�k�w_��mE���89e_���9
����ً+s��g�g��IB�6Sz=�%��#&�8BW7z�]�~<n�N�����֣�?�y�Ɲ��C:<N2vz��4Ň���>��ߍ��b���:�g~Jc@	���d/�I���Z�Z�%D���L�s6�s4^��@�J03���/:����^\<<��b������Ƶ� ��X�Y(_GyE[Jg�����|��c�`%~Ţ��/��!��t���4������O[�����X @�=�:��$BZg�1O�J��Ҋ/��_�2QA�W�G��e.#���v���ܰ� �/�BF�KxExF��F/d%`? Kd� �Zs��Z�gIp:�;wx��HKݒ�	m�}��tsz��:vӦ��e�??���`�Mw8�SR��f�k�h�
w:a���.��@����1\E1j���xl:�r�^�Z��͇Μ[�fI$��
��)#�χQ������Q\i!��9��0z���5	x��k���W1��:=�H��$l*E�����2ǚZE0=Ak��5 �"
���WSDc`g�x������^)z%�a�!E��f�����]ʦ����]z]��h�Qv)5�y}���I	˜�=���`s��դC�	7ˡT�ث�̛��Uy��o�������#d�:6?&����?P�;���ZTze+�iK�gş�Wx��vp�7����1�z	N��X�7Ġ�Ҫ����vx��8E�������>e����h��A�]���,k�{T��iaͩ*�E�d�Y����f'��0���#)<����Y=U-T+��)�� �V7hc���A�k]�9.-�D^�m�}O֣Ǒ8�Mb.qcv����
=��Q���8د���IɈ+#cS����{���o:�����6�:�$+Į�3�LOU��k�jN@���Lڎq/^u�@��+�����mֹ���Gv��]�|�,�mG���lWbfH׻k@w�uk���H�Y�yQ,��F�A��=��"����q�� yJ��L��q����53å^%�a.x�eIsS����%W4��%w��ߍ`(A��i�����"]��X9գ���ה6j�me�6E���<��������l5��AR�
�W��)UTZWrۅ���J]%��}sP�j�w���M'��'V۫�Am[�;�;K� ��-��4�m(f%$j��Sz��8�S�ժb��x�3�m̆>��U{R^j�%_X�uk�)#����eĪ��}�> �76l��׊���taacrɉn���"��m�S\�u#����t�-�O�����"�q�����_�#fFm<Qo=�p�����0��R�h�uX�f~�҅[wW��ɱ��a��ܦ�������^s��"b��W�;�NEf�.�B��y���^��û��T4��I�BxDp,ݳӋ�^i;� �,��|!�9��l�����d8���O�8�8W��tF��q6⡦ʴ؊G�H%V>��5HQ�x�,3C-�4��:���lABḵ���ቺ�P3���ԗ"[+��|�,ʭ]4��ذ�H��10<��Љ~�Wd�5'ѽ��X=@��\]�J	��L��uk/��6��>;�� L���og��V�!��U')
� ��AO�
���w�<f:BfF����a��#L�_��-�ľ�������V�C�6�V�$�C����
(t.��:����Ϥ���������~V��!n�#�	�j��#�@7=���1u��p��v��u�C�<���Bh ޗf.$^<��f�I�)�+A���
J��{��g�X_���̾wl���4l�̆H�SV��J�0X�d�Bh�u���y}�Ơ[� ��A�CT4��)7���� ����>���m��#A�	>�i����Z���m�qLa�_Kt�q�dNJ�O���p=�Y���_���#[����}�\t\3O��0E����4�A{O7��j�k�568�$����V�~���|�p�(�-�=��".���}�� Gs��ô�+k5�X��%k}����n�[J�˄�@�B��5��[��[Biu�(v:m����s_��3�!�>f/��\�Y O�Y�.��NX���U��b�$��o|Z��}*D�;��X�TQ��+(tT7q� �m����6ސzM��s#���f"~���?k[r$�U�հ��Oؒ��ՑpФ��g�R�׈8ʉ�|'�K���H��[G�"�e��;ƶO���Jra��~��y9|e�<��OYX���h�b�ӟ�DŻ޴�����]C�c����Q E����C����8;�5�VA�ه�@���U�Q<7���;Sr蓣cg7�*!]q�p���Զݗ:�r *��\���o���\&4��N^�bR�����Y�U�؜HpoV7
y	�8t�J6�Jڡ�M��|��i�����*��e�7�G����{)�P}��.�9g�vU}�sȅu~�����L�"�^�<fx���i�齆����!�����VDpX9x�&��U:z
�M|;�{���	n��t<3��XHG+s�<Q|�T�����/O�FY�-֭�쭾���+��Z�D��W�4��Y*s�l�BP��f���fw��(�X5�C��+(ě
�4��v5�@<��L>�pYŇ�6a%YK^��gť���?C׹K�V�2�۴�����rۑ�9�b���D�;}"p�D�t#"u�z_��ark�����_���	�9���M#.�,����8Mw���3�@2SB��+e�ua�
�Yy��;������8(m��Z	�D����O���j6�lȅ͹��\�U�z����`c�4A��2�AJ �4�x"�̿x��)�B划."�ؐ[��uT�Ak!|C��t�\�~�>އ�1�!���qC�L��~�-�O�
F ஶe}p,n{�Y�+���4�L��G��\�+4yQ�����������]�=Y�9!���`�ټƜ�����Fi�$�^�mw)���@���OG���k�t>�izYC����j�P�4"�p����+A�b[�����}��_��P���.�/u�_���~L"?s����̷]����>�Eؘ��hךE����,��I�ؗo!&�wDe\mk�Pl��:u����F<=ǳ�EM���ػ٘�F����M���Toα�z�;��률\��&��Νq�Z:m@�7�µf��V��;ٜW,�������}�~��Z�o
 JC�$rGeg:�b< ���r@L򶐢:[(�`Q9��0eք)^"Zfcn�Ӧ&S�80����5�g;��F��(�/,��K�G�Z��t�Ic�(v�o�5���Q���
y����틑if7[�'V�<�r�綘���M�X
�qP��~��ü:�R%yĀLQ��Ԕ`T{�;�7�%"�uAi1Q>5�_����q����%%�����d�l�sBMQ���~��}h6���-W������T?�o���+�ғ�
�!dޫ ���!*�~�j���������վ+����K\_������n�%H��o>ʤ2G~�@�
8�P��B�/���v��Hx����?p`�V�<%�3-I�f��f���/�
�-v8����w�=�怰Ɩ�3�N�Cw���ÈFƴ�H|ղ0���uV�"H��BFb�6#���{�F� �XY�w�MlZR�?9�o���u9J�y'΂�����%�
<��i����q���D� ��}៘s�2!�\��B���!¦}{�Mg�qX�9�I�91h�w��-�V���/�B�.� J �t���~4ABy��G�:���P��!�6T��ոؐG`���ǵ�q���X5�wu`�]��3�f�ŝ���~��aaV�s���O��-��4Yw�H$7���J�FQ�#3�r�h�ck�qt�G�����C�.{��5���-���Q�\Zi,H�����Ƃcb�����k�;zRq��n[�"=#N���$�EOoV�=p�NN>�
�^���ع���3�����M>]l�ܦ�ϖA��7E��K�:+��ʈ��H��G�!(���<������G�F�cF͐�i�UJ���K��y�K�0	���6M�]������m���C)��g��C�u�I&@檛	|���;S==7���݃�L|_���X�kz�3�C�f{��)�����n��t�[����	��H�n��a�5t��!N����~�4Ż=\��-J�i��f^|��R�_�JCZ��|�B\L����jb��p�2��w��κЪ;Dxvj�&�j���@�ԩ�]�'?[8��c� j{�a�9�S����纐��唊
�2�K�{��Զ,������y7�y��d?��؜:L���ҁ*U	�|Tę�8�)��@{��-.��|1��w��ܖ���^�a��Y#���i=�aoƋE�bN.7�r�c	I1�R���`�6&1-��w�΀�2�{q��nLqR�ȹÈ�����ZdU2�;����Pn�,r2	!���@>/�T|N�S����q��PT�����;�؁�q�6��(5��D٫���;B��	�� ,�+w��ˌ����
�eAI�o<fH�X�Q<a6m���E��]�H�XFʭU�̔��U�Ho(0��>�P,�]���Gʒ��۰�Ͻs�߰��P ����5J�LXLJ���`����,Ke���O�i�]�z�Q�>6,�Y���'ofS@8h��;]��V@l<m>V�C$���3�{����ۋV�~?Y1���tI�:7T�	�v���4���HN&�Ͳ���ay��lA�����,��v�myk��%Wd5^7�&,���u�� R]˙{u�?�����Rg�\\�W�Uq�tZ��\a�(��F�ݓ�{��F���9}]�Q,�����"��"]������20~�Ϫ�L�	�T'�y{z��U"����8���;��I/�pݯ���?�R��zp6F�~�.����'
7��umbe�E/]���"غ �9�����l�L���9��B��L�q
4�'�`q��Z���<��އ&��M�G��c\H��8�4�,l	��ϡ=��讲	K�.�W���_x?*���9��9r�H�ft��K�1�Vj��DQB��zQe�f�����'�d,����yda�w60ma�`'d�s�j����<\'����f/�Ol9��h�ǔpZ�a�зM��2��O��a�c��IB�4C�,���������ROK���U>;l:��V��\��H)�B���\�g ����PA�3�NHO���!�RM�� �Q�v��L��]d}�9$|7�����Y���sӔ$W������.�o�����4*��O<�Q �$��,���T9�r����`����]�G�w�����;d�n��M\�Pe�@Q�}iÞ$3��Q���<_T;Gz��ڥ��A�~
*oy��`����/Z.RV����zY����<G��A��\�jW�����e�R�d�����:�"�YNV[����|��*F.\~����gͧ<#~��:��Q�HU�BT�4������ux�қ����~jD�(7?#Y�ߍ>B�-���#�v�>0R6��TE+%�&��Q��Ϯ��UM55y{"+`�:C�k��^���U�I;�c���b�NԚ��apfգ��$[w��.�(���Y�N���թ� �x�mB��G�P�P�Q��e�c����������d��Һ���K��z�&�A��V�A�N���p�=��.��B��E��5��<���0����Ms�*��Q8�o�[i�Ll�d�2d���x���GI����8'�b�;����M�A�'�������4�h�^z�J{������d>.,�۰��"�`IP�R�$��<ͽy5+'&[w��#2�!�X�^���\���{��.�v7�v�wS���;C�"9����hD��F�-<���L�	<��{I�/L�VN�8}�l���F��_�|us������|�ưH�*�s=JYa�QV�~�u��b̤k�N1O�X���[S8���:yZ=��8<I4욢%k0l{�y�Q�=�\�c
m5M3cP42�CX��5����ˌ*��G�wQ�	�)0�O�-�B	EC����_�u�$e�<�0�ȹ���G ';!3j �VOQ���盽FZ]�|��$�B:��Ҋȏ�ު�9Ur�p{a�
=��C+<�#�iu��L�,�/ռ`��ER��>�z����IQd�S���Q�����rv'C^�����v���-c�>5���r�s_�㥮�ӝ�V���x�B#���P����G�䢶G��2ܣG�.A�G.lh�F٠~.�&�w'�����ݤ1hniX@�^�d�����޲�v��Kj���m�����Sp26[,�#�^V8nd�����lpsVC�B0\��_3|�Nݵ��e;&�mo�bs ��������H��s��g�z��É�?͛��v���bu���d1���Ǫ(�<!�G	�b
1�-]ӏm��n����n���Ta���&G��!�ԫ(��֟��݂߾�m�ƭ�
Y�Hk��ݎ��X���$���LU�58��U�9�5�"�zKFi;j��S�
��-�>6�k�KbG�f�~�� |��BŖ����5�w��+����',��I�- �h9 ��;�����t^A�l���)�� ǭ���X�Ǔ��sT̸�26�T�K k
��`*�q�v,�sƶT ځ)siޏ-�Vm����O
&���a�R�N8���W��b3�;��nM����V����6j��X���+=�즒�/�'�;&ZՔ�Τ�W�־*�/�F� �D�w� ㎬�����
ĉ� ���Q�84��wKa:>�c�L5�}uM\��R��}B�:<;f�l� �ψʘ�W����1}4���Gw� |�����\|W�s����'}���D��#1�~�M-?�x���s�BZI�@��O?����H=9`,�p#	��>�U)g�ť\���Kg��Q-$[��y�E4AcJ�� ӗ]s�(#�g����a'�HXlxVHYEB    73fd    1290��m�#��;��5/e)�M��1�?�=� �`J[P|h=ȂE��b��hE�͉k�ɗQ��X&Rz��FW�qG�y�܀�/�@PX6��7�V�P�悔�c���Ў �v�����n� �?	�o6C�Y�#P�Q#|�Z��x�W4�����U%�u�rU{	[��H ����ڲ�k�G�������F╔������Rޤę*�E�xl�q��j��pğ��8�6�S�_��N?)���� ��S��O4�rd��Ϫ�zsɗ��A�T�� E�.t{��J��s��������1ZQ7ƧR��$����q�÷�Y(`$�d�9E0�yF�-�S�o�u�.����%�Zr����DvLJ5P���!�ǲXU�8�7��y� ʼ&��6ǆ8Y���������8�bRtM�c��q�3#Qv���#/Q���L�����Ð��='w���)��/��t�i�2z6��L��)��>��ޤ���Wb�؊xd��H����9 �7~��vJt/i �@��g���3��8	Y9�t�p`�͑Ka��A5�u�����X$�&�s�+T���EɁ��1aM�"b���8�Dy(˫Պ�ϫ��x�L���2�KgtD���yH�=o�1�ݾ�BjrC<�Df=�a���8:�P�c�&��,$/f�i_/�~Ĥ��f��cGx�C~AR��k�捨�4�6�qi �M��,���(�V�!x<
�I������EՃ�0�o�;���Dkw� ~�C����p�;�$h&B�[/��{�	H�d���';	c�<F֙�{��p��uS^��I���YkX_�&��Qp�{����>5d������0���4�6;x�w��Hq�S�T��N�Y�/q	��f�T��h��s�]d��u�v�/K�D�x�4���K7��4S��R�4%ʫ:�3�(�n�!IP�V�X;�����|>̆S_�eǄ�'���	�\��כֿ`&�\����2m)�&ۤ�y�o�|��x�E�� ���+��Fu�`���]/G��1������n',���@A߅a_�C��C^R�#��4�N[	X�1����@4i5U��A;v2(�Y�F�r୞�b�bj����Q�����1��uV����1�_��Y��D��%1����Z�h,8Y�e����TG�e &�i����*i� ��j�c݆*���RVgx�S��0�a&�ie`��?��������g����R�ܯN�L���p���ڗ���X<�:�睼F��u	;�rô�\Y�'�ݖ�Ǆ1UX?Y]�z��j�γ3���:�n��-�w�@iM���	�j�(*ƵO�5	\cl�Ȓ$���7ʔ3�%
w(����jX�<��VI�L�
�śo��AO�8���VzE�1��2�]�t�S	
�k�����(��D<NO�PL�?�鞆�i�[
6*8.��$�Z�=7U��/d�R7�����bN��,���	�G�3N�3m����e�����x�ʇ����y3�	&
��+3��8G�@��K��pN����%cW�R�Um���"Ea.!��������no�\j=|t��._����S��J�/����v	ˏ�Ĩ�ѡ�@�褎�nl��U�L��.m$��xuOt�f1��EGflFRC����U��	[ېO:�¢�Y��׭�,m���v9A\q�0�ϡ��F5��1�Eq�u�u��SL@$��1�H��?3�5N'F�
��ё/I��\YNq�G���$J�i�N�.�#dY��9�~�i���w'sW��x�e��x����
9e���e-�%�56�Z~bO�y�:�oڠl��M"����B����`�����:}�|�ڛ�7��Z5\FDQ�Hp�۔�>�g�}!y(~*N��������:��E��ۨI���(Z�]F��.�b����5hj㨍A�v�ucm\;��Eൄ��a�冠mN�~��F���Rel����W<*���l��o_�ʋ��eg��&���${L�L�-i�q�rӯ�q�� o�g[Q�m"�oI�Gj��"g�����K���*�`��q�:'�(bS��"�\�!n�ќ/q
C�P	��f;+�<��Q�pت���I�O�;�v��h��F��G��DDo�����HPd�M-��ս^��p��e�'[`N.�K6��fj�i ���St�G��Ǐ?�c1��Rㅧ��O�T����te��>S�����B��c�6����Ib`�N�j)p;���,ׇ����a�5�Bv�<�n��/{~'(�����]	K�������� ��¹��2�]X��'-��$Ӓ�oF34�e��S9;�D�����U��+K�<�]���%Z�}��7�G-)�������i/rqu|��
f��Gt.>b����"vM;�5�զ�;��8�YS�Nٓ�}0�A�hB��N����hL��<��wB��al̬�A���޵��S�;T��]���'���WZ��\�-�w��F(�Ԅ`��?��v5W�O��o��u-]D�5WiZ0�I�LhGR��f����	ͬ
���[g3�udUv5���JF���3�������2���Ef����c��&�X"��|y��'^���F��!�*f��0�"�_	՛��IM(&о�$��/Ԩ=|��nsXi�oGHYf�AH*-g�rKp��`�ak�c����G�H��e�?�O��Z�Q�]X�Mv]���I�-� B��xi1��[`��N��F�y{�v՗�?sb[z�/��2!�8���X�c͙�d��nCK�Cp/S��M��e�8���أ#87��^��%ixEK�A�c�>�>0�ly�r��=�h�k+U�����zܙӭr4����[d�Ya�jS���
w]���ޥ�a> 7���G����C��l�n�VO�!&��2�T'�q�l0���ƽ���J%M	����Ĉ\�G�r��Ɗ���)c���Ê����C)�.����|�L�ݐ\�u��s���AH���|��ƽ�Ҳ^{��2�3����׺�fШ:��d<����442�o�aPR�:�ǖ]jH�h�.|��J����=�88�9�N^��@���7Y�Z�U��s��ěa�-�6|Ճɭ��Etҙ|��*J�Wh-���<'�ŋ�?�`��^���ǎ��0��	`3	э����3�z��T�� ���ѭD��!L�"ʲi�A�)]ɾO\��!��ި���{�̸�k|*U�F�P?.;W���瞻"i�݆�f
0���0�I����q"c���Yq-br��0n�r˵��C���0� ��Mnl�
�p_#^!s?d�'���J��?���Xr �X�u�ɩ1pQ��vě�2Sߎ��r���x�"��)�L���jG�$ ��6��2��N�����x��$���N�vj�ؠ(�?��t���n��dX��S��X{�������7�:�ϟ��v��z���w�ӰY�� �j��s�R�M�c��\�YKia���6,������匸� ��S9�{��e�XM���?��W� ǂ3(�>���k	s~¯*�"����s���E�"�$��g��K�NQ"d�J�o�.�1���2I,jH�^�k�L��3���i��m���mʙ�(�}T��k�\��E���Y�,�WԿY��H+H��ݡɃHe�����-�����
�1��Q �S�	�r�j��1Zm��}yaҁ�^r5���	�Oe��NoM=>�|F�P������A2�t���U�6���c�tn��5礕ɧ��+��
hEyx+�/�A}�������\�R�T#!<���璡�\0��9�/m4	<�^R���[9lnj���}��	�OLa!�����m]p�0��s�
bʕ�]�d���ã]��.x�.�:�8�V˴Kn�J<zVt �F�?�����Q�dZW��Z�l��1r�����LI�K#l�.��$fMn��Ge���[C�h�{��+���p,����x_ ��q�6C������^N�L����=W������xw��BU@�󄬁x'��h?��a� �@�iS�ueɄD�M�!w�2_%֊CB��M9�(e�&�(ă.�晫C���:�c�T{w��7V�i�8�M�0$�1��E�����+K�ԏ�/�sx�M���G��RF*�� ��������&�Nm�41�p��t�o�q8�C9I5��x���w%3Y���SF�!��<r�R�"��.}�05ަ��Z�6�A�c�u�=��(Q�d>�rH�xI�(��1����R�yO4�����Sźdi�M�ܸ��JZ_o���0#2G���v�di,[
�=V՞�5��
�rR�p���f�Y�����q{k��@�,:��Ժ��7B���7������3�[������Ή�_4�r�f�H��9�!�eջh��u˦���[�BV���	������,Z�d��a�G��WE�8�����y�wl�X�]�MD��g~��yt�)�PV�+S�$��T��!5K��󅟙��h9iH�ϛ� �Y ��8�fc#܎��b�n^��7����H4�f�P�0��/ې|.�^�y~K�įz��=E�;3K�eǂ��z $�	ꞅ��_`�K	\��Wv�I��܅B8\��|0�����r�3