XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{AO��3�/���������ſ�}���4�6�ƩK�ɐ�}Q��J�+�JA�]/U����d͝�������jB�P v*n~#������׷�!s�|<θ�8����kV�no�['R�r�F�=U��N�ǃ��kI��n��ꞿ��{�x�"����P&p�Z���~{\�����V����);�/��M?Ŋ�_ɐB��g'��%����o33��K]�{��(��T���_A����g7U��C������7�bڌy�Vr��%L�HjG!�_%��JO|��/'"V��QW#�*1M���D[�����a|5ޚ��Jc^!����T�p$^Y�*�E��沈�W�A��P�a�^��o7�>� �ÁSd	�o��K���6�՟��ǩț8�S�a�w��0��z�"WVe�����)mO�Kj�f��W�o���]Z�ţXu�*y�rq/���.v�a>szz��pE\|B�J&�H���éַ��8}�ܰ��aҔU���6o���:���C��Y�fۥ"�����N�������::�)�U���l�x��9�Nn��~v�y�'�tjy�H2T���HPK�"����ޒ�ǜ��X�������RU��&��F'���|��Ȭ��ڢ'l�*���������|��n��ǋkP��T@'I2� ΐ�ޯ�&\#�|V<��J�,�ue�`k%wf��{;�q�|>��!/��0J�Y-�z��o�%-��=� |F���7E��Ҟ;� _�6�����1|XlxVHYEB    f7fd    20a0M�g=�E�k����2{�/(8�6��~S��
, �*n^�`[�q9s/��Asb\R��\$����"�q�U׷`�F���ۭ�ΐ֚�}�6� �����������0 -�})�y~�O����ڃ��0�yީ��터F���H9,�&����Q�#�Y����f�(�ך�t��V3L���\4�tف~@Ԅ�<T�)"(aοXA!�|��Z[?o�[����0�N�΍�v?S.�CP"��zV��z-�'�ȏ��@�`��%,CY�vƓqJm�H|���V�K2���S���� u���\#+q�q�%j9����v������ ���z'��2ʶgH>y�Sw�nN�Y�۠� �Fp'`K���9Ka{E�@F����gc>�M�������_o	.N+���史���}��`8}�3E��b��4F'�pQ�~��������*���HO2a�%
���Gߵ;��_R�\5'� .�
�ē+�z������o��S���&�؃�p �:-x1Dd�ʜ~�gD���	Y�oM �E���.�3g>�}�@��f�Ż<�B:��D/}��G4��^��"��!��նUb�s�ݯ�Z{m��xP �E���B�f�'�=�}���^ir^2.]�m;�r�]�]���@/���* m�#� � ~P�=�0L<��P��+-�T�:�O�(Sv��Uc, ��f7;ܿv�l���9}z	ΰ�Z�\�GEɜx!�U�L�]�����k��.iP<��������:?>S�6.����=�k�CH]xr�6^ʚjf��̝[�_�����,�f�,���G��gAM�Si�<�Liڔ(=�;�/���^�z�S��A;��!^�2|Nw�����)a	ڌ�XC���:�m�:��F��ɞ�-5��43�3�a��{�׮Ӱ�@�s�z�kV�
{$iTz�%̩ ��	�D;{�~�@P
���A7��h1:#�jʶJ���טĚF�/;dZ (���NB؆Z�n��u��PQ7���(�Z�_Z�;-�(��<��?$�³Hcj7x0�e��y��J@O�A<D�+��4�	�6mʵn?� ߓK��T_����5��ҝ�eI��~試~��C,|�6U�21�C��Ƙ <�A��R��1��k�z4[��`���El���y,�ȟ8P ��zi�&̞_�羿eo7�g.�������M�D6�Q��3�z�����F��������m[||���,Ē�n쾾:�-��+j�����1z�hn��,��Q�I����`H�r���:�mz�0�Z�8���)�{۹�����&z.m�5M�����Z!�
^
�{�����^6p��rzf�B)u&��D�Y�s�Q���&����	�3v�����둭Hi"; U�-iFP��f�<V��0]O톗��1%q"��gwW�b�V��t��j�6�r,{��0R_x�=oL�6X*�@I�{�,-!Z�f'�ю:"���e�����a�
�x��o.4�]�s$'��Ѻ��\�0^0}�yp�K{c�/����������?��^�����)�)���@���tV�Ʉp7~�������\҅e9xK�?phKN�w'L���Jk_~�A�C��-��춵��\J���ߍ��=����-�4,�`%�Q�g
u'�	y5"�)������E�T$=�t�X�w1���PO;�y����wP6ͤ<_S�j�h�4���V
AI��q����c��Dؙo��Z�J�s'��t�H�=_w,u��͉���!���DlN�\eq�1�e�:9"�����)�O��deM8ҡ�"3GF��#;~PJg�N^�W��r�+�s<����T[%����Np&�wi�S�?9�8[ګ�Tn�L��?+���F/O*�:{S�m���-A|ܑ�-�q�\�M9~�r
&�Q���v�#�n"y#�n��;�����q+���a٬������13�;O Ç�A�}ם,��O�*�#����O���yL�1����8&�1�E�|R����2�ܫ���;�j�*���5�C���� �C��9�o(��#RH0_ u���5oEs�^�3��Ss,#Nٱ$k��	����w�"��?0)�^?�����W끽��s�5�{I����NN�:��Lz!C�������V�A�ʤ���<'��hH�S-ZxT]%]J�O��_��p��Q��-F�%����eI��=���?`��u]k(뤑FC������z?�6�P�"���Z
P&�L�BB���N"���R�A<���ږA�J�kI��g�on�L�����%/Y���3�;�zLo�w�~Ш#���T�[���
�Uv1��lQ#�\u��)x8�b���WT��hk����եZ�?O����St�L��62�W��#�HA,��+I�>%�L�P�h佂�7-�+��͕��VD��U�.�ū�x�b��ɣx*����E�A����r��H�|������K�P�I �a0:o=k)���>�$j��A����n	����+Yk
D�D���?�:���"����"���9���{�v@����t%�#?mUfl@�2q��s�Wd�H��F.?�1ɛp<��.���_L���E|���P��2ocA@ELq~�K���]���� ��([�E�7���nE�$����=��i��>�;)�k���U�f�+�Q1�W�#�:�*�ށ�d�Tl/Q��_m��c��ܝ��j8ls	!j���
ER�l�$V��o�Z�d�P�dR��G�ŏ�M�ٳ��S� �F�μ����<����6�i�V���/d�<�}Lh���r���oQ��΁�ѰZ��;��?pE$��,$\�9�����T��dxR�H��(�tV��^�O��(k��k��}�澴7�$c���C`�݋f����'^aۙ��R�^�n�J�&���9-$�zt6G6���H8���
o����Y��#�އ������c�#A����y�k�V%�M;W^L�w����G��k@esC�7��\G0\������}o��� Yh+���A��O������ˌ��љ�{VDV��sx�x��b�3P[�n�+:zl^�"��v���HCwO��=m:�ZO3U�l����6�Ԝ�"8紇:j����Ʀ���I��x�s1�KٜI+��4"����G`1�!�{(4:�ߐvVe���h �z�ʃHśC	6Y��������m彵�8Ԑ��I��z�ϼ�����
���s�#⨻�y�^�x�˦���U�p��G$�?�:zf�� U�'��k�:-6��@��0��nG&6��f��U�.4��	��]�P�����hW� ��ve{�b_�Vw�����"z)�·����]�8��u�e�qÙ��  ���q���[Ε�T0n�ʤ��1Q
+�yyjYh��)���\�4��&�q+�>�NǦ��fc]BU��Wc�[��w�q��u���G�
fqxe������&����m��:m}�I�jI���m�y���\�g�)4iR)dǖڬD�W�8:�ES��e�L�_��g����1"��H���
�FVJ�1l�% +��u�ג��ڏ��jgΠ��K+{G%�/q��#����79�1�0�ƴ�j�&��t*F�B�Hk�v�s��D��Ǥ׭�h'�N���l�Ր
��-7�P�?���s�Ȑ���=�Zb�yE͒+�T�#H�߁8pk5�c�k�K�j��s57,�z�Jt����6���L��ef�<"�5AU�cc��)�~I�.��C�ZRs�N���C�j��Ǯ=R:=�G̨����E扳|�sk�:���i�6�c�R�7�����OaVN�<NF�JmQ|K����⫸���b(Q��#Msxܟ���M�z��Z��=��n�k;��f���I���,�񦭋2w0l>��]g��j8ULx�M��ޥr�����XY�/W$��7��S"��]���G�3�ZdQ�j&B6��Xrf،�=��'ܽ-��Ygj�B��R�;Q�������~9V =p��;�&��Sc��������J�K�bO12�׼��@���m���������=�+����"��j9T@������SZ�����qf[�zZ�uYql� �^4�Ȣ5� �b#�p��
5��ZS8J���0#����q����H>3����������4 �E��{�۬U���44�<�GLV@��~�Ԭ:�~w�`[�S�X�-��u/Z�s~��"f�5���V�7��p�mc˩@����8�o���:&��O��2(!	)j_I�Q�B�9��|��{�
L��}��mg�
�ύ#�KX�����������9l{�� �������z�CC
���ceP�	�����HD϶�c�;�,���i� $�����^�'�X�U�����]�1�t5�n2�wG��̳��s�Kx1�d;�\���|о��x�nh$��U�V;�����h�4��s�	5��Ό��t��i���'$j��O���&��2����DWj��M�� �r���=�\�Iݹp7'y�J�i5Z�B���t3���Rx}��=�]9�k����hl��֟�[�#��O��������_��dUJ�(a��8ׄ�42d�N�8(;h�w�G�*ϸ/�4��P?(�1c���6#${�e´o��|-���������ER���X P�w��!3��o<�3C�/RiڙӾ�4�Ѓ�7J��r����		c��Ѱ��q\&|~�"������N��=a��u�j���:|6�p�%��*u�[�#]f��Y�w >7˷Z�����^b?�����١�Vyb|���4vk�	�;L� =�������I���FG~�\�{*ݥ�u���1��Q�g��^ҥ7va��(<���@*��l�ε���_���Z�Q`��`��i�ra�aEF�|�!����F���>6��g�#0\"E�:�N���X������\�}rɽ� JP�yt�s�I(b�o߆wm�/R�̷9`�:���TY�}>����r��c�p�bX�:$(6�PK#�8D?�l�w��
Qn�P.u���6�A0[Zq��(��EO���|M;��^�@�|�l�6r$��#�5�}:����?�Y&�k෣ V��nO��ec7f�.��ܮ'�?BP�]h��:�ĸ�j�4?A�3��y'�e[%*	|�<���#����ܮ6,������TW��E�I3�;Yy#�䅨:m|[}x����Hr74���������@5L�*R�w�d��vX\�2����\�^%�H��0��ǰb���Q����(��K|*zML���1�d�=�}s��oi�|��E*�N1r����q9Y*�bo����d����Y��M;��%�atD�^�ȏ�v���2W�U�,[�xp�-�j�Ji[��Uyr:�lOBw�o�����X��(,�	1���1t�0��<QcbJ�޽v��6�B���M!�T�r�2� C$.v��rd���c�����jm���!�����n)�T)|۫��(&{�ꙁ�Yӕh�M�u���4�.�p�z��"{3nR��MT��}P����ݮoT��=����z��lH�Th��Z[�3}�߈�v�&G�_m��@N|oWs���f��G���-q��8�oa��������RK{5������g;�9�����~C���9��M�Nd6=65);�ug~�C[n��i��8�,�8G��ǩ�"@,�����!?K�]�w6�)ݛ�;Y�d:��O�q��&���m"�D�qh1��	�p��^�cbPZrq(M����\������I�#
:��p�m%<6b�L�Y78�O�-![B]hC�?�F.[��HP�#2������Yd���t�D�n0��H�).��-�Z宀�&�+/;2�b8��;�ԥ����f�C1�ˑ��
LD�ct���r//aa��?-� q~ã�X@7����<oY�X�[�[��1)� D	�v8N=A�� -��o�3bC&V�����R�̒��U��ȯ�4v)���Ҵo��s�t)h~�t"���w6
�����F�/B?��T=�B* �́qӭP�.]w��n��dU��ƑR��A��sT�[�ν�BL��E�N}:�0��q��3,H/���L<Ѯ!���P��
���k�F���}{���kge:��f���YTi��ҁ�E0a��:��ɮ\�إ����@S�?.�;��_u[�]{\����Ul������w�%�*��FZ��K$z��c�卲%�.�e�����o������k�,�����p\b+����{1퓝�{9��W�F`I��Txڼ�jm��	LT|I �W�G��k���S4� Xe?A|T�M����4�2�2�x^��v��G��z,#�[[�{�*�2���h�u���v4���jQ���O��r�S����O��TVI+7�;.^�5�����SOh�~k39uNW1p���k��Y�HGmI���B�Ģ�ٚ�Rx����@u�Dj&�u�'|��H8)��],��S����I�6����,$�l-���I4���Cq7���%�j�����#SG��p��4�"����&��_X�KN.�߮��1,U�́�1Y��X���Y˼�/�#�Zw���Zx��:0��(��!����{�uMҕU��"=>s1�j@��v7�Gw��VP��׿8U�4hRWQ�Cͱ���ʂx�_�q}�� V�*��Vn��W�@acd�(���P�`5�\v�*�^����bk����������`Z,ŀ��-��$������˛��խJB.?�\�N$�D�?dk	���B���P�V(;���'
8����v�-��/}����:ex��B�� �LT��f]��P3�~h��Ϲ�Wò�E2Ez\Q��(ʂn�nD�EG��^�"�v�ΨPg�����n�BMr�.���Y�8�"��>+Є�IG�2��,D*jV�\��BDc��Ǔ��҄x�������đPT�7H?-�ڍ�]s��~�soq��� mbQ�H�[�M��eA�5j�ru����O+�l%
ӱ�F8 @�C�II��ƭ_Z�s�]��J�x���Xo-��
F�rt��!.>Y��0���3�ҙJg�=>�Ѷ��;Z�1�=��
�~�������I���F�J�ǌ�� �K��MD�ݾ��o�����0�̄�(*a�k�$�񊘚�a`q���f�\
1�w�ͫDC"������� ꤧ�^Q mD��3��2���loV-|y�D�#՞\�����fi���;z�v�	�uĢ��@z�渨�gQ���S��BB�;nE`%��f�v���L0w��~���%��Ã�-5�	tY�����E��Y����2�L�t^"�Z�2je�o!�*��H�bPƇUB���z��/�p-���T!:X�a�4iVBiC��[z�ZmQ&�;^2R��#:ik⪞q�wL�.�>M��6%c��,R �}\��bl�x]w,�|�~�JF���u�>p"��G/�f�9h�j�������w���nV���+��%��ĺ9܃o��}Tq��v�K)��\��8���g|�����xZ���L�/�R.<Xu��0B(���w�ܡD��2A|
#4�Z���]l�@���R�<4%JRZ'(0\�c���[g�3�=f�B�n��ȁ���K��4 &@��������yhs+�%���$W�ʸh��Y܋�Q<�r5La��ׇ-n�Z���'�����5[ܗ�u��iIcΤ�Vd�\k����|�}w�>��(5u-�H���2H��b�Q!�����¼�/N#Q�{ϣ8?��3Oegw�;�S� R�@̕fP%�]�xh�Nb��l]?�$����1�J�^U��o����G�C{K�x]���9@�E5�t�Cy3�y���Nn�$r�x��W�pPG��f��R�1�[��)x"��[�o��tb�ﲋ��t�zi(��& �4��m�&�򉕨G�0S��L:Y����t�ee��� �y
+^������:���4���ZӰwW`�w������!yР��Yì���۞�9I���(z_��s�7Solp�P�H�z��*����"+�K�'�tBh��6�H�Γ�+#��;���i���.WuL�׿$-����c5��[����Mg��"j