XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0��O��&�W�PX���~@p7
�$�� ��$}�ثN�xS��Ryn�B)���vR�����Smw/ʨ��xs����y�O�T3N��x��a����Z�p�E@���8f	���� �Q�����O0�D ��u���
�M�*��4^�^�T;ֆ����C�}�f*�7�Iք���N4B�����ݼ_X�.�o%u��Z�Ԉ<�ҝ��bo��E�����/���b����cl�f�	jm��5j���~T3�ۥF��E�*TV�=-o�'����Y�K�˖-F債�kJf*6"Z^��1u��ƉU���|�H������Ӫ��=�BOt��|�Xe�h�&�b�u-.ߩ;����`Ma�{I�3ko������Y~譀ik�v½; m��^b�<ZM���5��(=p�נcy<���q�����\��PE{~I{�* �{Ǿ��̰�����[N���N�vdp|�E{��n�2�T�q^s�4��zkH�5c�O,	���cs�"0�'O�Vz�5��} ���~U�$��rtlJ�A��3���+�VM�N��I�Z��4�@H�<W��)cl���1�lwo���`�Y�XE:�6
�i����sH��ϗ��YG�"�*�EVt�����B�k���_�f�^y\�Rs��LG��D�A�I��֯Q�D?�R�Kl�*����T��M[��l�_�w�T�yD��^LK�P�Z�s��=����'���!_dg�*Z������a�>���u�XlxVHYEB    3d61     ed0��k��X<�	�Ͷ��TR����^<����>r*��hU�8<HWx79������5�T�}���3F�EK�� �S�6\2��<AGR��V�kd]0&���q@��(xU�R)]�g	8�׃���|
���m���c5D�,3=�6�E>p���vs��h����C$)C�@B��웴�2�ȈD��ҍ�J.�'=$h�xP?�]�
�~[�r�w��u�/�;3�
Z<q����ƀ�0���%䶧��?���-z�!#Q��{P�t&aU�8l��IH�\�ѽ��ݶ��8"]��<*&�Ԉ8�
���w���&��8��C��@N|�d��/�#B�ZF�6.��N"o��;H	�]�O���\��"3Z^:�8ӂ$��҄W�G
8�moI\w�9�{$
c P~������B�o	�S\#SL��6����X|����UiT�Ȑȿw�a�z����6\�u҂���B1�hʭ(��u�O���x��v�o�V�oRb�d2�OǓ��FRT7�8���<��j�@�:�e�j���մ>�إO:��rL�m�E������]p���#�a�݁�!j1�5�Z��I���~�!��Qߎ>���W����n�Y�5�.O��p�``߈��J|���/T�a����6����)�U��W�1~V���ϔ;��t2�g��t�&�?�g���vT�u�tޙ��҉�H��C��z��t�����G�E͖����jb~d��԰�����k|���R:�f�LC�(�����^���9_e�c�}?q��������aW�_�l��
x R�g��]��,d����R$�F���p���q8���C,wM��NH��`���X?5ٙ	�b�����d����Z��puDj���Xɪ�]{^�n��>�ԝ����4�d�d�D:p�*�e�&@�,\t�&џ�Q�e�y��fN��"��t� ���b��O�{Xh�8��Q� ��v��޳4�j�BZ�v�56�q��5�OC喯�?69��K�Pf3 *�Kco�:�8�c5�o'�J4DEq%�Y�M�=`	[�d�p��l�w)*��=*S �+�rF��|]�{q�[H�K1�SȤ:CǴ<�k���R�~�@���<XL�����c��eI��rl�|u�n�k{��QA�/0���G���_���%��#�<29���!@�m����k��Kn�?g�p�������]?�L�	��n����$~����e�:��T&�*�B��wE4�h ��Iv���>X_.4/Yq����Dd��|��0Bf���9�Rrn��KuU%ů�/�𘵺Ћ 0���2�¢��k WxUE"A�i9ں�^��o������r*�;/����hK�rJ��y���v?{����^������2کnY���֛!���k��ycMh:����m��}����	�v45:��6vX	cP���6mBlcUsL��
z����6_t������,��zT�W���X�shE��/���I�{���}�+�����D=Y
�qP��)sCi;��������^y�?4�ujC� �(`�yoƪ�|�C(o���~�����ʷ̇��b@3�ʄ(����k!�9��R?k��92@v_���P��R8��+�JJ� �GPlPz�\'�ˁ��h��U�ɬ�����W�i�86�7���F-�ī4���L}і}��7(?���<j�.N��D�i�U��8�����~l��qaj��20�X1W̏K�\b�:�{(���;8�#e�Z�4;��]��%e@���L���y��<�a,�n�ڛ'�F���~g;���c�4L�k#F�W�<�g�n^چ�7�6��l0OG���"�3.��1�
kP�I���Ƴ,j�7�+	��QƷ�,�r�b}�F������Q"��bP�&�,�IA#`���81��n�A��T��,@�:����HV�����M����t��P�c#8�4�{��Cf~�3��`�ѓ� V<�>f��o+&�k�`�Asw"��z̪�~u��t�.r���[�M3�àE:�Z����A�����C�A#��)y'�n��>��Ha�ܣ/ѭ�@�1��O�yQ�3�T���������X���|g+��kGOW7-�J
��2fZ���[ ҁ�>�^t�p���L��fu������n$�\�,h����+��;�?o�7iyB�ʪH�33�(Zw6T/q���Bx��Ԏ{�I>V�DXC�
Z;�ڊ�����$�F���eUH�,͝��M���߮y_��vvf�
�V*>��E��n�ק�����cv�-��8"�R�N���\���e��H�˒*�Q��$�ڃ�xz�7h.t&�έ�Dƞ�JKP�4��/Ȳ�>�����/χ�A
>؈�}��V�^���,x������Ԕ�c�80LRH��	�@�q���sw�G���9�a�}���Z�:������Hx������.Y����*i��~�p9��()�F�f�a�>�2J&��Y|x�= ��[6vIF�ǈ�`uY�Vc�|h���bp�Svi��y}8��(��eG�x(6�TN�:�W����f�J,)d����M����$�g�G��;�\�'w���k�A��I�cd � sָ&�|��p�!�)�$؍!��$ �e���7XgkE���Ob�ֽ�4��3�<'gfYuce�;ħV����5�8ة�>V+���sl�.���-�2!<�u�o���������EeX:.� Iur�WG�1\2���^*�O��������!EkfI�&��~jm���	�`>2�3:� �oD�ԃ�J�)����)ý���P�mA_M�:Ԗ��;`6k�2�00@�cy�h�YoL�A7Ob��U#��1��n��m���BǮ#���WM�ms�O�cZr�d���.�z��e�S������9Q�39" �~���s�=�j�To�
�cI�~�ⓤy+����J�wJ�:�d%�{�u��6��[�Yf��26$z h�l�Bo?aO�Re�N��#u
�R�/���7
�o8*p��>��2gl��\��S��Ы��h6gŒ�b�B��f_4j{7-�n"��ȫ�h�`5���v��wo�N�k�_Dh��8K�*��c�����4@ޞ�Q@qj����B����ѫ�݉�
�;m��Je��l�I�[�ٕ�ɛ�뜏�I0`C��E�)�'�_�\H�w�e�?mB��b�%��bZ��3Z�7���o�%����S�����f^�kXA��&|�:g��F��]�`e2pR�x-���vM]A��WzkU�\k'��V��j�S�Z��/�}QX��+��QĬ-J�g��m��5��d0���Pd,��0a9+�$���P+bKN]��IC�]�7q���Ј6���[7x�<0���ףFE��;jPƯ�#�Fu@'ϼ�rC�)��r���]�9��R�A]��ց�
� p]��o�A����v�蟼ܮ�k�"�EqNڒ�&��}]�߯'�O����.�����jD0����$`��~~O
j�L��=\i��2(M88\�ϣCؓ�X�$��(q�O~����(P����'��Bg�{9�*/�����~��om##�����ի�dǡ�a-u6��a%���]73��v�h�~��"58RzƽH���Y��a���^��vm��R �I($:	���rY�c���[F���y����R��H�
p!