XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������:Ү�����;R��O
�M)s*2	w�*�����/�9�|�Ў����4�y� g3:|�:�(�٩ϴ�h�t�Svc(0�f<<���1`��P�:���]y�9��g̭*�ڱ�7�w[5�VΫ�
��PW����B��@��^ �"l���S�:�1�9C�o��T�(��k�4�H���ot4���
�eR�+*;#��L��.��LGETP��Y�d��S�ε+0���:�9o�z3�#�f��) ��W�D�x�ͧ� �s����PH&p�A}
I�F�z������C��}P�AB��R�[���K8�#��-��fS����� ������ ʎ4^�!7�P:�٩IΰG�`]�e�&+̧r�(
��o"�W�ZpXO�YuF2������J�a��c��h�2�t��� |��{����a��IP"�	��/N?�P/PbG��/u'��]�\M&����Ѕ���Ț�U<xsy�g�XT ?x��m� 5b���z'�9�V�ټnmZ%�k
�p�n�ˀR6d�넓�4/R��(r��1�<Nt��v	>����[���6��0����\�.r5���2���D-or9�:5.�������@ n�wS_�]�Q�3C��}���c�N)��9�&�-LJ���ji����.����O��a�d�-�r7���Й-�cwp��\X��`� \�Ͼ�(~�Q;�Y$�5͛~&�Dv�J��;P6|��iȜڞa-�x��M��v��u���&P#uXlxVHYEB    8990    1bc0��mÏ1�A��L�X����rA#40�?$�[G�o1��l�!��d�eU�4�}�g���g��{	c�5'����f�d��O�OE��V&ʬ�G�m��R�غ/a~c{*V�N7�ch�<G�����=�l7�/�4E�A?ڟ�����zt���Z���t=�ou���Z��M6P�{ ��L�h�N�D�����쬓DY8 ��(O�4ZŊ0�! WD��?�U�� ���{p|���+�W�![r'72�t����*Q$(��m�#
� �|��!ShO�}��� �o\*T%���j��N�J�(`�x���������:��ɍ�r����[M+�������bLk�/5?]`ėK��1��b�M�����Պ�NQХ|��� SgxoC�~~��
��%E�����i�8�^o�q�Z�7��c���珽�z�,�<H*A�F�.��'�щ��h�Q��,C��ѹ��eU�GS<�x@��կ���2��Ix����N�,���tڇ��=��g��^&ځ!���'��f��|d�!rT�����R����}�B��y�� ���z�e���*<�_�a#�̭?�qje��mo���L���h����(�T��s���@�V_E`�@,�
h1bҒ7��~�j����'Ӝo�� ���Q��[t��zɮ���Vk-Di�ޘ}�#7�D���l��cK�H ��K��v��'򢴼�o[S��gi�;���֞�G�G�˗+p�Ǡ�q
�8r�kj@�({�����{Κy�.��o1»��올�"�$a����8�a�a��5�K4/���[3����C��Q�/�̰w�������,�I�5jyZ�]�����3W2&F���a/X	���T�9����IT@}�L�U�uxzK]G����+�	�z`��#Z1B�����,%�:��F�m�%�D�.�ʲ����c_,Gh�L=	dpIe|�IA+`#�)�2z����s�V[�'Uq�41��V���{fr��kܴjh�: A�������������xŔ�?�/�п�:w�[!�R�^���zJ�O��
��]�AfC��J3�d�����SSBۻ�[��������b%���!���\|m3�ՖYCy��`q��8�|��Ŭ#�<�R�|� �A<ߴ�!����'���	���@��\RhM�u�6sFV�V�}y�Д���"���#ժz�~��_7�:_�L�ފ'[���?L嫿�xn(?u�XZ��J�+�P7�ǁ�$}��������$���a�jLT�|��p꧸�_���M^�7�8�j@y��ʑ����Ĕ�5��Y��:�TyX��.Ũg:�ǛF�?c!��Z�8џtn@Bdl_��m�x����7��9y���J
[��3������(WC,�/z�,�A�����;�+Ȑ��Cp�~�:_}��Ë�v;��ȝ*RҦ��`S�W���1��ϭ�<Ҝ�������[Z\�sJ,�L���k�OV��Ғ�
������x��a��)%"N�բ�=Ի�ΩŘ��nI�W�ǭV*Urc�"Ǯ%�T��ʑ�8�b��`�*n�.�Z�1�B�G����R���u����6���C��Ź�_5��	,�.�B��C�ժ�Cv��VX�w�C�Kz� ��[�{�c2$�V\�b����+�A�X����L9Q�Ц ����d�뙴����9|�����=�jyUW�U��36���D�M/K�W���)<�h�����[�#��I�0$��S�˺���X}i�!�I��R���ex��"'���5n��&�-@�4���PF��VYY����)�/�˚��u�'��:�$�?i���XW�m���L��$��,��� b��iW��[�'�햛%6���i��I��tό�~�o�R�U��:(���߿e�M�N�y��"ȋ�Fyr8�50���p��l�B�+L}�S�9.�o��6�!������\`��2�1\ה��La;�uNO�[�4�5s����I�7�w��4�Bw��]���	���f��8�^�v�-�|�6�W �z�}p�OZa?���"K���`�U�E�#��l��#�~Rqw�(��|fo�&C�ԓȵQ�ܙp�d���H̯il�m\Ȳl@��P�AL�y� )=Ơf@3���J�8�. ���l��Q�z��y�@P�,�I
M�  �]�x{6�S�Vd[�6�Y�5����j����=ϩRuF���'�N�k������tj��aZ�mB:jUZ�w,�T��W�b&��<a[ 6��&���[���� <�֌*�0��Po�����%. _nWz�!�E.��	.]FFzx��`M�O�J�� 1l)����G�}�]4}�������o�9o�;�dX.zwxYUCuG�^��L���f�<�(紗�Zf+w:�Xׇ�x�i�e�f
+s��i1�z�Ԕj���V1�]�1���7Z�K4j.�����N����:�^�j7�/�˹��c��yѽ�7H����KiFK,��:��HE�+�^Iǳq�W�����oB/Z�l�W�Hu�|K��r&ϵZ-+K;����¯F~Q��;[���򝷏8I�r5YI+C�|��]H�Tm��u_�f��˥L���3q��~,�2�õ'����"�mp�(I�EWWQ��œ����(�M���Pw�?�+o7�!aC#��`�NV�Ŋ�E�P2V�+�08x��e��d�>�Scgd�����v�U�-�K���j<�QF�X*�
O,�-vŏ�}�IYO�*���l�g��ֶ�F�Z��#d������ �3�r��X������J�jX�ń����P��P���B�ر�]����I�(�����o��O���e%z�A	�uG*�x��
W�]����*��ctx,?�0�k��P*��G�-.x�¬o��d�#���H�GT�ƑW����or#`jiT桫��PU^@kO@-!SS&�[ɨ^�{��[�OmBaƹvJ��|��x�6=�C(}��!�I��p���
+�Js�hR���o��+����l;�N>�7؇���Ҍ)�l�LeC�<�z��\�y�0Z@)60�	�#����}6���� �E
�.��K=��(\ț3�@P�[;xSDg�0#��R�O2�-���V!*!4�X��E1:��m�u���.����l�H�y"�$V_F:2���oF�
l��E#����;�>������4�>��>2$��Ň�Q�[f����/Ƈ�q���/�W�Ͱ�
$@���\���j��0R�6�_��A6 �휋Ws� �l�HF�icǡ�W���S���h���د�=aG� ��/����J\�{�Յ�tbF�W�\�͍����L�C�����:qJ�M$��lKIJ`P~�����l���u������pDȟ������/��E`;��N���'���J�~�I�t�њ��ǀ�1_LFE�&j߅M��ex�6s�W�9*�����$�':>myZǕ�Q���A���^#x��Q{-�P�<�b�`D���YjK�������lP��Y����Y�i�#�;F��On�eN��3?�=�6i=C��mT���U���`,P���+Q7|�c(=�t*L2�F�>�]��3O$z#�������F.b�)����)�*c�l����M�����>�'���?�\�Dd��!�9�̻UZ��)J�x5y��+x5̧�ÿ�z �B���A��	�������A�OT�P~Eg%�jY�d�n���"(�&~�
�v[���[6G;
�fg`/k�yu�sBZͲK_cK��a��;�I����B���h
�����u��@-n{ʜ�W^0�����R�p��-{_��׀��H��dǑ��{����p�z������V^D]3��	��V:�g��(]7��,�C+���^4=��&Uk7\=�e�W���b(c��7�~6~�n�ϹR?-^���b�� B�
���+>[��I�c �oe��*�%
��~r$s���j��z@"&�8�6�n��V����-��}�#.!�����(��I�]0���,�[Y�4� �����6���U�ԑ��y5^嗒-gS�S ��9 [ڠa�\N�iZ>����-c��{U��LwR�\-��y�&g _0�]V�S)�y���Zr��b~yF�������h�'��E�b���6�/�o�k�="W�V3������Q���.�k�/�%X�YVƬ)��O��%��z�z9��]71OJ�W�9�}$E����V%����w��9�q�Bܝ�}���R�a]��9�-���4�v64p'pb������O`[E�>�چ�dN��������6p��K:*!�"�G��������p2�����@N�@��q)����L1ą;*�!9y���S�O�L6Y�& ��+
�d�E&˓Ү�����N�=�l��(��� z	7�d��VK����o?��;>6���G��W�q�	���Mo�#�Օ��%�GV�+��ɟ1Yz'�'�
X̾*��� �R�ƚ��[�q��3k)T�� kL6����S�c��+�"��8r]|�mP�2��v����c�oPE�)kO�k�v}��g!�����.mH��i�	��$�@a�;�9��*�ǵ ��6�)����ȶ��6(ZU��3X	iW�}�1�>�g�vD?,7�hJe��� �#þǤ+��\�*�~��.c��z�5���< ��+�?���O�_Ġ�zt������/��cF�����X{G�����xAGAiS'm6쒈S�L���u�Y��<�NOQ�.�K]?��>���ZG�SF.���5IQ��?hͬ���UD������������1O�JVC߭�ѥ%y�(۪�gA�>�K���*kl,�M���,�ǜw�%<��E��y<�,�Z���X��E~�S�ބ���
���ލw���\�ɯ�#$k��0�f�Ձ�.nt߯6G��p�զ�D9আ�?��ߢ��p+9�9T�آ:�Sa�&�@�hZb}��sŮc�E�j�)c���1)���oL�+�޵�H�ُq(��-z7�!!�����y�X��۵j�<i��x�:�~T��Z�װ�3�^ٍ>���\�'�̞U��,��j.��[~!h�}t��x�϶\�>Q!�?u�f�E�&f	j�x(�Y��O��c:b����+���K��h�?f%�1�Ý� B��y�|��QQ'��t��>�}�����6O��|�����z̊"6k�<eR�g����1����d])ď���┲��י	�]>v�,5;8�5\����Y�Q�w�K6������3	��@���;(�4y�2Ɵ�@>�i�
�=�	;���I�뀢����yDm[=�E����ſ�p�*�%���j+�R۰Me[�ʣ{���;��ze�j���
����	)	�c�<c���w��4��uJc���涣[��.��pľ��V�;��D�|�xթ�'G��Y:W�}�cC|��]����H>�*��C�/کf? ��y�b��#e�blmx�£%\���6��W�?�Ͳ����C�W������c&�n���i�:8x����?	i�U;�p�'���T��F���Л���G����qq��0���2�9�3o�ܲ�����(�ˡ��l�p�i�W~����7uM.�'f����7@0�sR^� ����o�$���%ȷl��Y�FG,CIO$x�1ڱ���&݉c�p�M��ۿ��f(
��'v�г���x�� �-s�m.�MbQnN)���|@�sT3}UҴ��ͯbDq�{��1řUJ�lt�:| ��l�G%�������AHf `�k��r�(�ށB�_�ުe����iAF�����*�c»�����Q���,�)�
rn�_�,��fk�./�N���D����;��BV����a���H��gL�}r���;���6JU��sl&��:G �Z��c���㓟r����B�Ε��kח�2e$�M q���h�$ؖ�j�]z��Ӿ�_Ǹ|cJ��T�mfՕ���*T��`�3�I'���K�_�:�!�J�/2��gR�+d.J����y!/ڊ��?���Z�����U-b�HvT��YC�)"'S��^t�>sx��0�>M���N�P��nyӹ�o����Z�.���8�Xb�e
����ֽ�����)�P�2�Ck Q�W������\W��E",��(�{.�Se~#�3}1g�]O�/�b�9b��V]�/�j����>�-IkD�)���"�l�V \�U��Gz�q��P<v�,k*��Mw+�\�R�u�g�@��J�X�*��<��5H�����ߴ��p�}�.A??��
F)�
�+:oi���`t�������H�3�,� �:���E�Pt�)V����<?|jǂ���lw�0���3"$]���/�`���]��'�U)��X
n4�|{�3\)��L�n,����RZ��uK� 2��.�<�]�F2�a1!����|�yz��j_����*r��-��@�ո�X��k�&}9/;M��E��b'�L����^t����h�LX�����zC�µ��������RvL��J�)�Qj�t����zjP�$�T��j`we0t)�B�^|S��.p�Bbh���GV�g�ƹ%Ȁ��;ř��5���Y���t�U���gz�l�����P/�Ȅ�Z72�lK(h�ė�c.�Xj� :�υj^_�+\�a������f�Z��c�a3�^�;�]�nW8���l34��,q��j�M�@H�.�L~�G�"�5"�k�9�ؕH/��߆�]�RQ��#2;D���$�,��4fV�?F�K�0��ko�tkb;g̏��ߊ���N<+��E��c����H�����q=5�WcJ�O��$̌�mϋcE�?���6��2�M<�5��$���фN���_��0(�=���9�G�#M��f������ǜ�Y[8���������