XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"�َ334���#W�|<�����ph8���ு���ۧ���4˥ �F�����*�W?�#[�*FA`u���7|��N�GzoQVǨ���������|�i�j�Y��Y7X��1ǉ\J�Ȱ�V"6K�PC�&�%ſY]���p�R!�T�!�����t�Vl!��c�0d52�0M���<m�����;>%K��?V.PM_�?���[`��ކ���/�rekb%��z�#��*u�n�����J���,&~ے�E���uv?� �·���$�������F��t^'�l=���dC)v��2޵��V/�:�b�}�C6����;=w��l`�x?�Z`�h\�D$�&i/ח�/����Cݫ�,�-�>������,Y�2O�����r2H�ԖԖ<�ig�4�w�a{P T�fi��}o������jպK��6ӹ�$s�gQFJ�fp	�&r�q�í��|c��H�8��shȽVkI�]�P��a1A��BpX &���b��������O�/�_\����LI'�&��# ����=��5ϛ�-�f���3`�HV��Q>���-r�7�F[��Mȁ���5Sl�ߋ�v"�L��8Rn���9e���?��V1�1��u@#P&���ލ�S�p�-^�<���*3��$�&ɲW$H+F��7�xWΑ��nn��DS/�o> 0��?��A�>\�&�S��K�c� ��M��z呟A��o�?jB	[��ײU���pf!P�d�)'l�X-�,�l�>�f#�h��qB���XlxVHYEB    6534    1400G�1��m3���g�.�I��hџ\ƴN�J4�p�}6l�] ���8�X%%79vo�:(>��a�f�7�䪀�"6�������0R���S��C�����\q�}=���X�Q�\�]�b��E� ��<D��m��I��`�����m���{���
JM��wS�Hv9��e��h�|f�����Z�k�me�j}F�^��Ȉt�)����;G����G͗+��1�:	<�Z����3���� �|�������\�t~�<A0�YK��Њ{�?�F)D�Ϋ w�~E���X���>Du�'�9|�S\	�	I����!&��q"tG޹v�PZw��i�6��OY�3�gk��(�%�9p `,3��������ª�E�Ǥk� ��Ǭj��Rp,���%k�L+�?QOuPڴ�7P�}�=��~� ����ҟ��\o{��bF�	��б��Y�&��y����O����O)�i+Jt��^�]���d�G@_�����9�!_��'�Η&/ĭ�I[��k%W1����z���955��2[���f��ƂGv�n"�� ^�����{\���|�vޗ��HY�~��jA��>��)ݏ5�Ӟ͹0!�4O� �j��E9�������E1�Z�Rޘ �/�p��t��&#���j��|�h11z�i���a��O��U�(�o�
Q}��)��J�Ϙ,�<mm7���<Kb��݈�v�`�>~e�!;�]qf�ڄ�^��]T�."�F!ęy�R�_bà�������trb�3��_0V�����A}��k�G)���l �}p��fZ�-�����[���K�WpK�m�怘'�<��q9�M��r`�7��m�e��2W���T�+����~hB�����Q�g��n����׍��H��%׺#x��SV�K�� �a��c:L�������$T�� z���C.��ǒ[0<Nu��Y��R|����l6���|������<v8�z�� K�q
�X���i�����cT�X�#��=�J�a:���> >)�3G�
�����i�5t	ot�Q[S�8]�ZW �G.��׿�˲�,�7g��'.M�#רZ�
+�Q82�Je�^Nk ۮ�:˯���=��oR�q{��#��`������@�e��+8���B5g��xW9��=ݢ���^�{��	b�1H�a(��K�[3a령 �`��5�0�?e��t��0={�R \���[dhw�;�Պ�֮n [���ou����Y�0^~h���}_��ٮ�A�O[+N .<��.�C���:�Z�� �?4[<�U���L�E����֞4M1��ϫ28�B
�)���e#�2m0�^66f��|~�P�����j6g @�-�'�����Yc�Haz�7�}�UЙ{�r�u��|t��T.Sv��=�%x��v�����
�kr���5�:OӔc������FU�>=�'
�Fg~|!�4��Wy�w��cJ"���fo��u��������10�ʶ�}|ȷ��[���S[&�������b?����c�ްjvKƧ�m+��&	J�g����ٺ�ՃZ��rM�O{��Y���:�n�����N�t��X����f��
�U�^�<�r��ўp#R���s��T������<y,fAy���np�du5rgb��}��T����J�h�����uvW�7��H�����+ӢJ�Q�{�dq��|G8/�fH,W>��S0�I�|'��w�$�,��/b�t�HO�c(7h)>T��6�T����{�*��h$�$1}Q���{í�	`ƀ�[�{�y�W:��L�}��4p�v=tO@̳N/��0."��1Ul�۩��b��X
 �t;�f�E�ϹC�� .������+���z��QĲOI�]�F�0#UE_����^�
|>w���b��D����:W_���{޽��b�5Ho�.fW7u�O�i�Oz"�o���^�� �62� ��/��������LAn�O�N���}Q�w���(=�ězh>]�����{%7�K��%�޺9?�����Ȯ�l���BEu��Q�����>S�9��8ǁv��/�G���������g
���u�p���9)IL\ ���X'��Y��aE�0J'�ê�_yP����BY*�ÂѰhJVqgbrsYZ����7����di�����On>!��d־��Y��Z�z��<���2.�P�0-�Y����n�)�&��W[F�͌$�,���:�$~�c����Y�������ag�IW�&!��z ϟ���2�Fd$�#�`\H���7�7G55��q� �ঢ়�ׅЉx%/){�G����+tu���_i<{үMh�H�U��fBo����F�\����Si���M�Ѡ��:p�q�
{��ӓW'�$\ρ�?t�[iQI��£D�,�uM��X�0O�Vxx����C
�R��[�6�!UghM��,���Wt�u���TWΠ�"��&T��8����~�a��c@3�
)�ǉ�`#��k~̢�%�tB�\���'�VJ�!��r_����Gā��9}�"F��7,UV#z��W3V|�,Rz>�e4��OdR&nGW-��BW/ a���#&3`�����Ԃ>I��7����G,L�s����Tm�_�1GH,�T�P��*(W��=�H�P��#��#c9��,l7���QO��y*ٙ�iB���PV6��t;[sgu��H�sJf���*1k�%7z���&�@#�8d��j��"sm�.�R�(�s��;-�q���AG����-��l����v��"~=R��E���V��G�JQդC�U����S�>���Bc��.G jIz��}%U��X�G�@�>���	�	������v���4DHK�Iz�-�[m�����M
���2�R�? �`��z�6>��,`�eL��{�aD����>� x*.p�2�G;��_�����V~���3��t�1O��-F�E�˅0n�+�R��k��dr�U��<r��t�����,/:�Hu(8N�d�7e��H�Ԧo"{>�l�Ց�2�k�.��H�Ǝ�^��޲�62�i����ٝ�8�LUk�+\ �<�?Y2��>wGY�M�鮮��&uԭic�c�/�:�㡗n_}� �8d\�̟M,=^�I�u@%��M�!J�*��=
�1P���)o.k�~x�e�!��:�t��+��	${j�RjL�$�I9��u��8~��CH���(�T!�����b�JI�mŊ�P�B���K:3��]QZ6}�Q	c+#�x�p�����{\K 'F*~^�.�,��iq	�v<,0;���e+��_&?��@\b���w?A��RN�`�-�[�|��eދ�U61E��o����ɷb/�n�$��$ts�ܭ�*|�]5�G�>�UB�٠I��{�<�I� ���C��_w�Mڷ^/��"��{��
:7������%T�B<m�>B=O�]�ע>`k�`u��#
pO�$�-F�'����8G�{)�O�x\WM�����.Nx��ClQBg��Ymz����l����m���	t>a�W���*U���!8&w�$;6TH y>��ǡM����y�|��VBq)��Sro(��E�?�8��ˑ�le)���Yă�m����ki#�K�&�h������k�٘O����9����*qw�t8ki)T� =?`Z�V�pd-8A+�uy�]�7 3.�� �sص�����+3��U�Eɞg񼘽��]&a��-Z���ם��8�',<�����4�4w;hV��!7Q�L4�N=�-���f�!���w�����r���}T���&�����] �]X5st����v��(����$�fd*ph�.Y�`�7���U��b5j]�P����)2m���Gs�MN���/O�F-^�BR���8��I��#�<Q#J������Ş��P8tr��}��3)�=lJ6�O�ۘa�g���K#����u��<�P����o�Qy���I+����[�����B�2i >b�=¤���/�_FG�v�*1�U����?�aIf��,#|�����~U�>�b1pjP���))��_ e�%a�ϋ��q�����D^�6����1]����/e�i�-;�vߦ
�sqt�	;Q=��~���u��-g�뷸
�	Ӝ�`mɐB@��d��
��F��\��.��"��!fR"�9~�D|T�n���ˊu����n:�2��֎���[/+�TM~Q���#[n��d�M����hGZ���#*��2d�e������z�M"Lδꔀ0���@�y	O���\���&�I7�2ռ�u����$�������Z��	[��������΄���g��Kς~(˿C%� D�\��U\�y&�(z�ߩ?*�$�|E<掅k���C��Z�<�Ȇ|_戣���%Z�o�cY�Q��e�s�5;_j[\s~��ɇߐ��l�ڂ�t��*:՞�L�� S�QI�=��ӏ�E`�W� !�R6��Qԟ3��~͔�ŐL��u�X�u�wqb���4��"9��e���l��,�FBYB�9|Fp�w�#olص�3�1}�qK�<0�w| "ߊ������r��7y��+i��J|c�n�w�u6�����냙�!�X���d�����]6�f�J�u6`p�"=� 5֖���\mg��/�'�M�;=�����z�w��\�%��B�c񤑬C��eڡ�0ơ~��� 1�0t�D�����E��������^��+$I�N�ƅ�U���l����<�7��	��@�K�*P��%�3�۪R�'�#`"������~B���@@�3{����T�U?6�+`dc+����ӗ���=�x�Yy���u�ZQiP+�����S/��V<wٲ�|�f��6@i>a���@�w���X|�Y�ǐ��IQ���N(4����
�R?�\7�հ��+]ȧ�E���+AM����Si�E �)���x�9@����9� ��8#�؁�u��Kv���ϏFF