XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���.�4n~boO�O�߄C���n�ٿ��P^��e-J������7�j�Ȱ;����ӹ��*
R�H`�!�G���b�t\(���l�g�痎��=�bG�/�s�a��#����O�&G��N���g���M����R@�+1;��F��lt�C��
J��*��]�'v;��H��
���b$+�֓�F���--������~Iu����[���N�B(��q���}g��O��!Šً�!S�΋x[�)�]�!O �FI^�:i1٣���E�;=xC����e�D�b�E� ��/�����l��D�����e���B�!C���#MAޢ��g�7����U���I�+ɟ��g�L�h��r�L��q�;��JQ����+ch���!i�=�ƪ¾qB&p˔`(�e$_),���py�,*4�&V�,��� l!��'Ɏ�_��,��?|x���,��cI�;e/ϼQ�l�%�EM�2i�+���$,�Ɲg�]
��JD2S`��������:W��W�ʽ*�_��U�(���C�=���gl�dc�E��
q�+�t���{��0�Ŧ��O3����նI��J&������BDL�I����v	JLPo��!^\F:�Zf&�+�}Dph��8iEf��x}�y�n�*�A).۾�d�+���P݅ƣ���.�	[���_'�������^���<�G]���̌R��Yo%N.�o�=��[��_�CT6����t���WXlxVHYEB    2bb9     ad0��H�*���4hrC~��`���5���hx�|�J5�#� ��j�'��,`}�#��皝����*����Eh*��O&}��:ʽ̎Vc;A����2}v7�`�,�y}r`����;a�'#}�kkr�eh��DE�f��]�e�C~��-K84��e��[���%k�q��TC#��W�Q�tɞ��)��U7 &�%�9v;!5W����ޱhK�,�߭i�L�fdi���.��V�3��陰�EB�L<V��9�ZV
N�5�C{,{(��0z휊�����1���*S햂���	*j���	��� �"߈�Q�\Z���ʎrщp�.�t_�����q6e�0���~��jxR�h�S���4��3��΃�o^��-eu�yElo�}�ٌ���ͿB�7��V��.!zp5*���ߦ��_��Rj�����Ǚ<��R�R���M;�`�����"��A���/8&��N�0ty��b��`��A��u�z�I���c��SCz�� ��F0?��9a��<�(�pU<�/�Q�C��12��YowA'�1�5ݪ��`>|
�1�T���E�On��hq�ٯ[]���o����ЕG:T����\��_����je��&�Qm�G����$�(�6	K��ϩ�������<�v���z�u�HF>,a^�VF��'�nzp�1ƭ�qU��^<�"?�98C�_b����)2&��˘:7�˓a4��5rc^ė��%Ω�`	\�/������Vr/�Nqui�������"�8�ʝj�}�s����ܹ�l	�9�8Hz�����Y��ղE~���Z�i��-:JF>�&Z�XF�8�w��C�|Uz�!��-�!��E�8�NˈI�-��yz?�X�%��B|&�_�m�ֶwy7)��Ϻ����mIJ��"1�ǌ̨�����{
���C���{@��P٭(DG=��e8-a  pnFg+*jm-�zkCe�X�6��������5Vg���T��p%;^
S}��4Q!T��gl7JnB�>-�����38"�5���D�t�n������2B'C^]�֐�� 
�����7���캅� ����;�[����&035�M��)��9���x(0!����X/���?6^�v"��k��>����;�}q6}(R<ĺ�I%:�Ҟ� �B��yEp��z6Fu�xZݢ��RYY�OJ�崺����-9i���1z���q�Ƴ��HeKyK���?oH����QgH�ѲX4����u�HYإW���f�p�l1��J�H/hc�����D������t`��%�pC~�P(5V}���\n���u'�\{��s�����&i1��K�ǽS��}J���[>�v����-fX�L���/{��&ĩt�������?�����Ya��?��?F��,�h�i��}�굽��������6�B�ґqFʩ�|իq@����Br-���t��W���v���� r"�o�����F�/8N��V6욏�r3|whP���lD����H�t.���,0�]z��cP��;tl`S��	��P!�RF4�����Ll�L3�4�g���\#P�l��7ilj�g>�]`;�q����[H�_s��#s1�_u��:4��������C;9D7C/���`��zi�6q9a�%�rb�x��Y�<X����V�6���8�J�~�n��JTi4'`�)���z�}*��E���Q�{zD&'y.J���Q�g� J��)?����#e�[<��+�iq4��?Q��Kp]Ƿ��g
�;�Ƞ.��S��VB��{Zr�6��ђzq�� X��?�@��ԓ�mi�y-ۺy@J����
�=r����jy޷�IEZ�=� _���ln�k�S>�!Tک����<���½+����I��0�Bh�@od���_2c>
��?�;�;�FZYK��+�f��1*.���_�����V� F��C߆�7#L����
xf����׫�ɤtz��P�0ͤ���ٲ;�=ix�Cz	-~q�*���葄Q��V�~~�?�MAf�K��1���t��{H��vx��X�$��ښ1!��q|8�"fm��� ���qA1gX9>�j)���M�Q]��3�eAc���1c-��q����F���
-^ނ�����Dh��4����<�<ȧC��=���f�����zM�i���m�d7))É�.�E�~�sT1��pbmM�����ze{�=n0;z6v���+��B�����c?�zq�rrȭ�<�ڿ��`��<�y�P��1��y�vfS�;IBE{:�t���y|F�ּ��FiU��G�@��9�9L?�FB�K#���Q3��h426+ �������V%�N�����s�n��]��Sn`h��]�<����g�2��ϣ��K��(�$%Ȑ�Ԧ��g��8a��������?�
�iZ�f��r+�g�[�j�31$�|���Sv*�0c�'�R�rtP�?��P�ּ��ڔ�-܄ � Q'Q�o�{Z�KwɎ	�v���Y��Ա�� 鞏}�=o�Pt�Å7�,rO&o�sh���	���<R��c�DLpv�^�,aFt����
�Fh"��VP~��K�.o1e�|ɇ��ie���b3�Eu��.��?DtrSy��G�ͦ���|��/b�8��op񞮲�+=qNfٳ��CW-U+��K5�Y�R��̜|�6y�ZQ)�s��B*-