XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Q�.��o����vo��|�7=�y��С�=�7"A����"��3C�FVpf�&��a琯��������4�
��V�s������#�k��W�t*����X��B��ܕŪ2T�o�0\cS3�^�ѫ�V,Vа2Ft1�7�~�l�p��B��۰4�� ���t�|�ӱ+��d��%;�1
΍MC����i����؁�~~��		8��}]���ˌ䩕���D������L��ZU�_��L��F��Ȭ�1}��~�ɣYy{�Iw��MZ@Gl<9�|�Y�|h����ls��]tz�<�c����(2~�O ��%tu�Q�/J����T��"A��<��=�Ԇ)m��h�:}`_��T�&��.��A�*���U�a�5��K�$��lN"L�#��whʏ$צw\c  ���VN����ȃ�Ķ��X��������ӯCtV�c�=�4�k���f��-�O���ƭA��3
/sF$b�S�QP�+/9k7#��iH�-H@�
ToC��ؖv��ȴ&�L��Ց�c$m���z,�d-���ސ1H֩:�,>܎�R}"g��^��G�[K_�+��F.�<�y5X�� _WvF�� ��f��g��R��8��>�&j���{�"O�<r��.ol�$ }�Ru��+�&���ѮgG������WV�\ĕ<i�H�n�52��up��V rٟP�t5�� �5o�I�۔c�q�4��҈axY���E��q�^r-�^*)��g�� �ʨZ�N�1��$��XlxVHYEB    1ffe     9b0A�OS "N�6d�Di��a��J��{d*4� ��<�4 ��A��#K�/�Յ�..�i/Y����y�i &y���3а	ڸ�Db��|�ѨRX��G��`;�d�X�d�1۞1����>q<�.��Q1���Z+Po�O�E���3Q ������p}3�ݴ��Z��#<����u�az���!(�Tk���k��6����P��-���L�����������n�T,�%Q誚W(-G�ʒ��i�WH�"y�r�)9 �g���/.+`�f����K]S0��V@^�X)�}DR��Y��\@:�x���L�͖���u}mlzo-s)%ިH6�f?V�.7�,p���ÿ�yu��֒����U ��i�S�F�-.r�W����|(62�9�T.�q"�hY��HҸU8��5?��2�r�r���f�� t�H���2�	���K��"�oT=��U���r���Ƶ����T���jx�T���GwT���F��h��<�m��ԻBٹ.p����9Ix�h>Ǻ�S�uN�̕q��l�(�3j����dvD�0�m��}��Wj�%�͸�2��誇��5..��SrD�xI ��qH��@�b��i�3�,0�U�q=� Z��L\f���(�q�I��>�;���ſ�P�!I|���͔N����Q8y{����5���tǻ��t�D[��!�$n�����+J0���n7x���(��ӗ�5�}����w��eY�1��
3?g�Ԍ��AY].�DҬ�<��)\��ƻ��:��D"V㕺#���{�>զ�s��*ޜU�j����c�!���Vr29)~0���Y�'�p�K����6 C�o��a�������+�����ɿ�ph
�O�����	�_�B;=�Q�ּ��G{�:��a�:�=�����H������y���e�R�|+����N�u��d�t������ɢ�lF^�Ub��RhōD��ޱĩ�����#���S�!�Xv1�����hV!��j`� 8�"��foٲ�s�h���"�2ۙd�:��2h��PE��|]����L�9,��Y<�!�K�ʶ�~�H��(s#�G�$�p
%�Z]�.y�s�����忒r�M��C�ṯ5�[Q�˃+-���/p��e�´m�i�yk��������!C�trHNi�x�b��)�CS�Ӽ��ۜu;�b�A��8��>F�:��?��dKyp�����[�\�:�T���N�]z�B��~���m~r'\MP#J��Z��d~��boŊiTg�_/L��W(��G�S*���U�a�I����`��_-�.�����1�*�g[/_�x��&�~}�15�<�&�9?��.`��Y���6�byϻR� ���t����?�K�e�;!��Enq���鳶F,��Ir�uݬ�0�@,]�x<(X��}�'fA�P�7�����NgE�V�)i�FH�D�V�	ݑ��M7���3���}n�s�DJ������5I�p��?����)�X	�>�Vʗ�A���tm��@�i6D5��D��.��uD+rӨ�&l���6�5��}�C�F�u}�� �+G&]�J��"�fj�C�$�ŝ�y���v	�p�?(��7�����7
%����j���x�~�� �
M�z�J�#j�t+�}~�O��������0�5����ed�r��a��
0a(��P����fo�c�����cC?���q+t�9N���2F(F@� ��E�ʷ����a�\<�.��c���yY&o�~���C�b��[��u�6�3 )��?��K��%���Q��Ӫ�|�s@���2m��&?��)?���p8�*�.���ɾ���=�-��6���`�l�=��6�bTxD7�\p�F
�=#���Z��6Q>���lq�=װX������+��r������A �m��k��d\�3��e����E��dh���b�(�bz�[� �} z�X��#0S�犞6��v�`�MIp�e�J�xEC�=�0�2�rx�4DF��rՌ!]�u}�a1E 1���$��{I����UR穉44���Ur�e��l*o�ق	^�)����=����gR�1��ϝlG)���Q8�ލ���>��~S�*���0�N���|Dͬa�#|���C�)�fԌ�뇄��]��Xa�7>�5��#K�� ���z�C�[�}_��,z�\A&�PR�7b�o���e�#��W�Z�:{�e.p4E�7��{��k r%>Hҕ�)����cx�8��Z������)zc;Y�	�nـ`@}g�}����<Mq��k<�h�j�����
F������`��"����	�F��		<I����b�^.��m�;���(y�L���/�!Ϥ��IyS�{ơ4yaGb >�1�R�ޗ���y�n~���R$ _F�1�T,������`���.�8WdN�#�