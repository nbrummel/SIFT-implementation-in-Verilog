XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Lbn�t&�O(��Y��1�YW4%K~��L�{A�(Sp=�Z�N�,�$�Y/��|�*�%f�	��y>աt�wp1=�:{$��
����5߽��]���?a����<B����I5���r�	Nn��p%W'$wJ9���}���f\�\��(-��ݾ��	��� �o�	Q����3��o7�Y���p�����ӣm��uKi�b�Y�S�}n�@�U��sA���^X�b#���@��n9��Y$b'�d�i�[��~���2Xmn�T��`��8���nD�^��㢃�(�hQ�d�r|�OF�T��Ӫ �[%V��I���?��O'�=@vH ?,�%�;<�!�i	0�m�$�l���&.:������+!
�'���@�#�Ssx2��,��b��s2-���;���a�+�b�JJ�����(`Ѝd$�V�<�0�����Q#���� ��jYV��.1���;�j�'Dj<�����Ln�u���tj�\��C
GS_ؓ��O9I����NtR)�f�YT!tY�4Y��<v
��E����(���֙O"�L���V�ѨQ�"ߪ�x�B���� Z��R2���d4�3���H�C,��(��ab��Ӛ��ISnQ���04F��&`n?ҋ���o��ͼ]�eU�d��7m?"Ab�-,\�Z�7u ��}I;"���	��VlG� ������7��MHb�t�� ���K_lgv�@;цL�K8ﬕ*_8�_X��v�I_�nq�O��1���6�$YB.�� Dj���XlxVHYEB    da14    2390g��9>�t��s��/���@)+VF���9�ǒ*�?�s�Fմ���KHQJ$B����{ba�z�����	2Y�!0ΏW��ю��L���������qQ�ۥԵIw>H��h�(�@j��+��kl��9z��[G!v3�qu 
���`���f���]1�-�~�Нz;��'�����w:s�r�>���+���T��$V*7^�&O�9Sd�{ߐ�h�|X��h�	ʨ)�ɥ�Bg}j(A�#�녪��%J�7���d��e���ƅI���r�6 ǃF�NTW<��ۣ�Q���!`(�� 2MRe����t���z��I������z���L[ޒ���J�Q�T@�T�t7(�V{�t%�GGS3F;�ViS�B� ���k9����e�7�Z����%AΔ�8+*Ԫ�}ko�9
2����/�lZT��U4�2~����Ir�N��_�E�ӈ
����%8�.���m]� ��|���Yݘ"�]E���v�������V�D�����t)L�R�ugV�z@U=�\h[�7$s���Ta�W�@����B)y�sS��,�A���i{X�z*9�Zc/
P%t�q�44���'�+W���Wz�����]���U�\��Hw�=ؓ�(�z!�B���M+��P)�%�Oa�SRH���8U��A>h�6ƷA'�$f�3��/Ԙ�?؃����hl9�u�R�nQ#(�>�}RTm�Kax�����{z�T�_IM���Q-�*>�.��I��Y��7e)�Xa�x>�|!9s�Od�6�Xk{'��[)_�B̨���|�K��,�!���&���`�W+ē��(�����.$�j�1��
M�iP^��D�\�X�e�⠅(BL�R����nS�a�����[TjD�|o�VRJ4�-��{��C㯖�ͮ��cɲ�`p"��D*k�Dt��#�K�¥u��E��2=�Q~����O��Q#F�@LO\ Y�j�Y9�&��s֮@����Ӡ��5����r�i�E�(�ב��]��H���t��K�j��)�
/�/���;��4�b-P�N>��~^�Y��,WM�+<�?�W��*��5�S<�w��g�θaTSU�G!���%�Cޏݥ�m�58��]<M��h�k7����x�ظ㱬�%���Ɯ)�M�i�wj�R�����Xl�aC�9�\{K�td
>�8b���BaB,�	�{��MH[g.G��&�)ڐ��i�n��]�{��՟H��t�C39PTTh�y���=�>�n�CG�lTHŢ��b���g�E���{�@���(���y�T���]Buj!w��������O�bA���'c�ʹ����|F|M�b�����e�V'6�7���@��|(�P�8�Dk��T�A�������qm4��](��_^�@,��twFB=�\+�ql����c����jaܶ�OsI����}a��m�cT���Y�aXJar۵�d"5-J]a� �(>Z�/r�^ÿ[�tע�8m�W�=q��0ݙ�*t���+ �N6��G/
����r|2�n��h,�󆎑_�fo����k*�2�f�]@Ԫ��u`��q���p�]�u9o��� ��#=nF�M��t�q&c�?�^�ʩt�f-�QM"qIc#h���[<�����숉�aa�H�������vf2�}��W҇�d0T��`�����`��"�wyE�"�jaU�4j�����9S��+�!�͸���/T6ߋ���ba�L���2�֚���ʸz-��=e�=uQV��t�œ��~�l�\��;��r #��'�ǜꆗ��~3�*V)g���4�	E�W����E�K�-~�P^��wd�k�����M��C�*�W��C���\��Ĩ(2�S���[���+j'��_)7��FvR��ߦHs,��4�`5f}8 ����Q���%�4��� ��fm�;�%�k,�Cv���T�2�}8U�!�!@o��G �xؓ����9�+h���d���2�-�-�u��ȴ���}*Jڤ�R\ ��x���O���BW���É�	�BTNn�!��}E�v�v� W�1�^{G��x��\kxXQ�j?!"f���<a���l����.���3B�l�d/���!:R�c�0d�D<u<3x��VC|���%�������P'�l����S��GbP�l�B�f�³�X�%��a�<}��@*<��������tHڠ��o`���������N�߭�T��s�0^w7qe jC{b��3]�Z]��(��?�:�0�d&��N�l�'�6</�����8�8�w+��H���~�yv�/�I��MY`�J�.��$b&+��.aÃ�Cn<��t�r���$êim�,�4�E�?�+.���E8CI^!�х����̳���'X���D�ʅ8�`��q�,Ka
�w�k���$HD-Yu}*Z	�Z���[K�|ҍ�FBU_~���g�d��s��f`{U���/���d���������6C�����Kx�(�I+
��K�CE�ݚ�W��/L�6�F����E�Fi�r<z��M�xnn�O�I����c�[�E2%f�H�R]$�OñխN}���!�Ӝ�Nv�x�S�㳮t0��tm�Ĥ@>��`0%9I�R:��G�z�m%�%��G���1M�eol��7�fq�V}.�`�<���r�T)��o���j��{��� 
����I�EL�tS�^m�_g�d�,��y��+f�n�u�Y˩����6��x�����5<���,�oH-���+a�o�_ƌ���x��-�;J� 35�� n0�
���iHRS0������[}^�ء�c�qVF���N���P��.�{�3��;�N���-��;?D<�IUyɴ��RI���Eaxl��V幓�J�J�:.�|�/����t;�.�.����l��2� ����iPN�C+�0\�Ǭ��'�+�Ƽ�ۖ��7VL|���� �q)��U��<k��/,{h��`�G�&0�3�>�]Nl��(�{�&�9�D��B����O��
+���BD���Ǟ���I�3�KS���DG�
D� ���v�4�Ő �*��& ���vṛ9��OT��.�U����~�|���M3/r�ȟ�,1}�F�l��~py��0��ݴ����[`�˗�}JR(�^��c>�
�K���]����������Ш6B;��\	�n+�����g��p�u�:�����"/�V���]�b�&�{��W��y���Bȧ��r�ɫc`��5��j'd�T[���y�(���zt0�?�:.�,�]����)�үr�^�V\q�+(�-�љ:��HXs�\���3�]b4Տ#�ئ!Gх���U��3&���McE���e��zzwI{��	eF'���tv^7qح�\3��ס���4"K�C׬��}�����M�&޼^�!#kf���\�yf=�ѐN߸\aڣ�k_i�O����wI�f�HZz7p�;�@��M.ǈ�:�1_��E�}xG>�2fb���p������X@"&Du]�G�.h"	R����
!��mn	�!EPT��|��~�y�$�_v�/-��2��;&	:1%�|L�T��u���xݨl��T�05s��a5ТA=��ƺ�g���&4��q��R�6�����4Q�������!�p
���nNSAՑB<PF��Eօ-X�U��D�fJ|��^k{u�<��j_G ?��~M�A���㛷-.�-6o�����n�����kQ%>�!��H`�Sj$I�[������1Np9�%9��N?H]Z�r$�I�)�� =�����y_�8����b5O��6�����ޣ�.@7r�+�����f��rW���N�&�ӽ[��'��!&*A�J��ߘ$���b���O�C���=<��`j�Ū0N�;��>=�ݤ���1��~b���\���3��8a���-�&�����$�;hئ��I]��ԥ��Om�l1Q���Ƅ*���P�� KᑮQ\Vk�LxZ��4�-�Rj�9�C����lP�_-����ja��� �9��c�H�9,ґ4�wܩ8�l:Q����ŵ��l�J��o������o��.�XD�(}��k�p3��r1W�B���e��>*�����x�y���;���K�-����.��3�T������N����n����_¾,������6�yk(�-,�k5��P<F��5�7�-J�P>��+�hm:�<��Gf��/	�:ֽڈ��h6b��^�ꀼ�:�"�C�{b����O�gӂ'�)�
uT>���~�W��Z���C�J�H{Z�h-�g�<k�t�*1O��\����gX��U�L�����6����yvQM)��&�&��xR�Gx�q�,�4@��QEnBP$h�Xi����{����a�ҘH�?Q����'�����Wk����Ӈ��O]���l������pt͵ŃF'��_�C��f2Hra���&E�[]Y�V�[x�#q��[��#AԌ(��id�/��#�.5���6�\�mO�q5�,d���a��d��F:ǠS�N�Ԕ���K��I�9s�Hh �ƤT?�T���X���M�̝��dz4=����Z�r�W�t����/Mx���\}��_gCD�����O����H�+o�|���(�`������j� �\�R�ۤ��}��|��j�C�F�Ӡ��@r�0�e��3=�b��.iO����[l�֩���C)�N��WGQDdje��9���~{����"���?����.���z�Ѧ$a_,����K��z���)� ��Bs	��[����Y,���%� �'뚻����N�h3]AE{C7Ӹ�I=%� J��8����/�d ��
�8���4��|�������ј���Zȯ�@��P��0��I�K^����;2\`�Vsb�=�o`�P�pU=�Ԋ�?Q
�&>��3�u�	�4?�5�\o/!h���{��0f��4� �EF߇�����}.�X��̓ۢ��:L����۷�HdU��]��*AOJ.RL&�W��Z�G܋���&7� e����Ϥ����7���b�U�KX�Z��^O�-8i>áx֥�� ��R`t�����Õ)��,��} �hA�k��_).ʔwJ(5EO��<˲=hy�g�W�����"�K�NnPQ�0*����q���}W4��w�:���������w�r���8�\�X�!TN�\���0꿆J"���X�������jNS��9�=���������{jW�ʘ�P��!fa,��F���Ai�H/�^�n����m1�ܳ�T���3"NBٮ����ːwr8�t�la[�ƁP��H�
iDͳ	�e��5`h#�����.�F}Oj8H���79b+U(t���>�ܔ��.�.o�<�^x�$�H��,rR�2֟=��r\�[yQ���n^ӭe8���)t�59ܣ,�v%3����fx��c��oU�#!����g��=�֕ɚ��޸/Ê܁�+��B� ����A��B��Tо'����M�i���^B�+�S�#-
�@�yY�4,\S,f6��U�i��2C�0�
��Vۼ�Ҕ]�.TǱ���B��j�*=p�6����X4�r�֟�9����`��?:$t���Ya*�t�M��K+v�����xt�#FE���Jo�DEs��:`�'X�./7�`x�`�8��r��6S�	��4����LbC��0����O�AYڇ!�K�����R�k��`����Q�_�j�������zEmD������|��j%��"�Z�b���=-O�L=fV��eݚ������ ���)V~8t5ԪKDd�v.���������n�j.�e�� %~a=1P�X+�3�SA{�G֕���OE@����eh�@�=EE���S��5�"�t�E���f�FG�5r��J������"�T�6{���-����K����rh	&�F'�
Ea1�p��n�.?�l0>����W;���V��(+���[����gm}��9=� a��N��θU&�5����X��WQB��s��ͨ��c�^O�d���p^�����t
���	S��4���?J�6/Oe�6�CS���8��I7���8�b��N^|��N�=��ԇ���e~����ɒ�=�[���GX$��z�AٺJ[e@Bj��b��ړ�ֆ�L{�w�7xJѯ)]P9Yk>G�^��[/��[��ZWoj<�P����P�ꌃ�g��L����D�Ph������|Fɢ�?-���[�7���s�:4<�!N� y�Y)�1U�G�%k��E��]BR��X[ڽ���-�zV�o��7��s͂\����9�G-�ty!���	rA���M�?
r��j)w,�ng&�XG��4��?ߖ.���(+C� ��}<��e�<�Y��I�����D��4��Qw�MQ���lޥ����ۨ=V�TP��:��ՃW�Uwmͨ������J�:��eI�C����~�F��8���v<��*M������@i����{
��C��i��3�6�)x�F�)Xϡ�k	W<���3%z5Ў���{�|�/�ľ�l��F�bu-|��]Я���J#�G�C]��1
=�9�T���~�)�y�{�ʫ�����������z����غ����Ic5aZL]Ė6��|V�k��['�D�}�&#OIY/�Y�44P���B0d���.$�U�xu��`������!d�[6R�Okb���R�s�	-w��rD=W9�*c���ϯg�1�!.܋r�F&��)XIlQoj�l�|+�G�q��si�B����RE�:M�N!3������͡�K��h�T��������3H`�W�+�S��=�AA҉''����XƊz:#�rij,`� 5�����Y�s�[c `Z���@��S}�JZ�v���q=�O����� {�B���fx����gh�[����&2;6��h�ha��E������:1��Z��(xIbR��~���< A�I"���aV�FD!���W}z�=Љ
=rδS}��dʬl��W�����6`BD�Q�?]!T ���F�F�Z~X��u��z-�����[���!:%�xT��#s��(7c����#��z�V��D�d &{�f+�=qj�!m`J&�w�~���Hh`j�����:q�=0$L��p�W40�^�_�}c9їdF�˴�R�hڿ|��k o���@���U�(ɟ�D�{ڲV�~(�'YQ�ΞI�˧��+.v��1+���N�m�鬬�ֵ�ȼhuP�?�ъ4ˈ-E��agg�l�C<%Єz2�d���`�۫�_�/J���������{ͫ�/�qH��)�cR�ð�_���2L�(����'���F�ϒn�z�{�qa����6&$X,�+ھ}�0y� ]�0��$�i cٍ��f�� .�H����>~^C���SO	m�)06�D�����-+���~�n-��G�gA�x�Դ�x�6���`|i�]�!-�,�t�(Xֹ��\�r(} V�d���e��NR���P�u�$̏.���xl�(��]��öG��Q8���D�c�W�EӉeɐ���¹�����^p�Ϗ��Q�,�xA����� nߓ�>њ@ ���lMP�G��Ϊ�fT���������ۖA��co2�ϔ�v"3l�[�`	��Rƶ����L8a��4x�7��t�8Kq�愶T��#me�Zߢ�-z �R<d��T9��eH�"�s4��ھ*��k �2��Q������wk¥��H/��C*��P�aS��@ǔŸ�0�eP�y��H����o�;�y�_�%O&�R_]֛�;��[Nv��&q�a�rm��{�x�Z����?ɭ�#�^/X�`\��Ȧ<>Qø-�c
e
������N��i�K-ss���O	���ŵ��E����Ȣ��J�9s^���Mٓ[�2�Q���&y�OzD��Elw�����i�D_ٖy1;Vo�lG�PC�ɦ(7hMpR�p�����d���5��U[c�%a�O)�Q�i*j��*�Y�\J<?�P�>����E��ΎJ�Հ:�48�j�-$4���h�:qڼ�Q��sʁ 3ewf�_��q�-,λ��V6����=�� �Ns��clR_��ڬn�=�"���c�u�0J�*zk�Ht`��u��$\�jE� ���w0/���A���6s6!�suTjD�\�6�.��`�<UB+��%�����=2��u�-ߗ�9]ngz+�WO��VTz�b���j��|)�xI+��P������;�%�w�C�G�O�x�T�a�1�+Ĉ��qa��hm�w"ѩZ�qʟΫ1���wQ��?k�J���Z�1J.���m�?4�9��̾��M�Eu�rn䧌���!����qۺ�S���<]�c�
Oeۍ|�6**$�Sx]���i��d\O�;�3�������{%H�a�8��Ǖ���$®(�4��3�XV\�������s��>�B����(��!̉��J/�ir���	����f��s7$M��"& �M<
g�5Ο�
�q�
Aq��[U�����店tj�$3��0�z;����r��˝�+��]S���l�h ��f�@ /ޞi�SV��Gg豪4n�z���eO�V�Ñ�.`q*t<�R�V�43�,��0��1�Z�Hy7<��9�l�H�5!0j��3a��ȹ;1'�jr b;,'�w��y�
������i���sxF��l�o|�\����@�b���Q�0$�0:P �����Âu�=.�p>c5[�~I�`@P&O[~�v�	T;����'a���Ҭ������߷�_���d�����4�h8d֖�Wș���!��	��;���YER�&�HE��t�k���eDE��͐j�&Wv>�x����>�w�w�z�$F�Y2=��k�*{b��6;(ٍ'