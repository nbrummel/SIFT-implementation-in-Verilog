XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����S�)F5��Wc����ai�K�z�^)�$}����BX�C�%�	NF��!b�EWѽ��Wr�EԮMV��Jv�3��ٍ�1z��ϴ��nK�����\!�u7R�k.+01L�"��9i[x.8�;���P)����`���?�,;0�U�ސE�1��5��5����V*�7��<a���z빎�mvL��I�^�J��'������@���»�o8K/�闀&��`s��j_Ⱦ��<�jx�#%Ԓ��s��}�%{t���7���h��4�{+�r�ap��و*+�%��IN+�>ku(�G/��pހ^�K�Dh`IJ������*4�x�_�q�=D�y�U���sn#�j�U�6.˶��@<�egǀOy�ۚ�m�����fh=VǼ�f�S
����s���9G'��=�6���l��	�s����,��Q|�u���
��6�6���/��b���SS��+/ogk����[R��㓥`�!�֟\�S�ED��:�$����ۢUP��*MT'9��U���9ܴ�8<K������TZ���A���H�u�uh�$=�-��Jp0��Փ�����1�2{5G��K���p��ժ�+u������O�=�c95���,n��i�%B��zt�	m�'�vf��-��&/(C��RPI��2��ڱ������#�Y�
�E��i� v��[�l���d� D���o�:��wv�]?�3;��C�0ޔaJ�.P�L�Zf:-��/:��;6#0��XlxVHYEB    fa00    2d70�%�
�)�M�X�sG/�jR����^��,u�y�ˮ��Nū���)\���L����J��yg�u�=[����'O�*�������4����T���n�u�#䥀��0n}\AN]@l#P�e�+M+�>�W���+�k�Uز�ߡ#Y!�c�/�|<���xP�yHr�C���0�߯�v�!�6�3 ���!"`	i�n�?�|Gan�뗘;|�9[C�x���/=#��8��R��=ݍ����F�"��g)6yga�m���,�S�����&�j�����a�^G��Y�}��ʲBz�KN~�ed�/��횺���*m��O^�T:U��o�a��ӶE���>ZɁ��W��G]���j�@�%eG{�wǼ,p����:�#f]y��sY���4�v�)�oqGT�L�մ��]���>th�g�Jp�9�'��rD�ihW�b1�"5��C�ٗ�Q�c7�S���7����>�S�
}u]���]Q�Dp�����u��c���u��������^��'��N'�1�Y"���MF���?v��8��$0� i"i�����R�8%�����gӅ�/��a���H���ϔ@۲?�џV*A�C��� >?f7Y�d�s�7����@�pV���;���K�F��ф�E��5ϥ�r�C���)i���$�c��;���ų�]f'��g�#�u�l�W9�HA�E��:�����Yv1;]?s��}g��u���$�4�+9�}�����P��ȨLS���� ��o��M*��b�2.�����		�o�|x�0H�J<AMp{�tΌJ��>���K&�q��vC?��)����dHxX��am���=/�T-P��{� �w�}���Y�:�pn���$i¡/�?@J�q��Gn��dr�qnT�Q�|�
�E��-ˑe�yk�/��m�u-K.ĉ�0�n��ή̣�NiQ���<#V���&�cw��VZ~��c�I�mdH�ŀV5�ydhq�������g����ƥ�&�1�=qnE��,��_d���h�ߙ����BG=�����-������+��0w�0����*�-P@}����/�=[X�p�Yz����Ha���+�c�s�J��hN,g���7[�߶2���v+�ab��3���p{��K|���=$���,E
l�g�I�'�0������,�F�kL�X.��@���K9��D'<T ���ƙ�<s�НTE^a�4���@E*bz�צhp>��%[����8Y�,g�W�$�.u��� G�ˉcצ�*iʽ�\n3oS��K3X�vGҵQ�̪���������ݪ�6����iR2��k"r3c���t)����ȴ:�Г�t:�i��ˋ�Ќ���:I��� ��>���|H��Ւ孢h��H[�#"���b��:/P�{QY`]Id�U�6�;��SB�f�,(}��
l���'�)�u&�֘_�<g��R���|�Uf�*0�kcZ��E/�<�|�L^��@��eN�Rl�P<*۾��e����E���he��EA�:c��O�b�S��L��H��oL���Ǎv����oJ�W5�C���Ӿs�!�2kE�+��[����Nŀ��=��^�n8�����a��6�n���\k�:�ݰ��<In���b��ؖ����P�\���.KO�S��S&��?TFH�;�d�(� Mp�v'/>�v��lL��R#_� >/��LL#�QOxn��T�;3�j�s�L19�7ܢ[Jg�%�@Mi��Vt��۹q�1"�C0"���h�������ubd�@��WJ5��/g�� ��W�<����%=�uA�D�M��[x�M�S���f��,��I���_}�*4S�SA�<���/��*u�K$�Kdy�����|�������P�gb�5���pOc���/��C��*�oj4�S�_��*k*�koSm�C�����	;����A�B4���|��s�j�Sj��M.B�2�~�tӆ��1��N�|��-H�6Q96E4-KS���6o���\�ڛ���l��E�9 -�S�V�H�/����F�HD�-jk�}�"��>$�0ԞgZ�g�9D����E����uI2��#�}���2 +�
͘�}A�A���ȗ���q4ַ{�t���������Q�P����b�FusM�b;^N���?�#с�^�-7>IY!�ӿ�@���uy[�WI�>�2���_}a�J6!8wwb�������v��e�O�l��0�^:9X�%���p�w��%�=�z ���^o:p�?/�%�k`e] ��0�$xnPE���N����|���r�5���FZ���������晵q��:8���;`ݗu�7�h��Y,�/}�{��C�����ck�69fȚ�J)���#���y
Fh���PK�"�n�� �`.���u�v>���q9�3�25bp���d˳����$�L/�s�c����DkQ!�&ڍ�{c����t*�;���~�h�ׄG�!���z�chX����3'i�BI��ƢT�z>�`�p��aܖ����	�<� <+:y�T�����Y���v"+�&�׈��m���{r�os�����B"!f�D�Dx�An*��م
$���z�6�-ac�P�`S��G,�� �(��ZT$-�E35��������p��M�O8љ��J��2"-#���w����c a������S^[5�`�	T{���a0oK2~pE����m%��]�G�5�kv/p�\lp�od>*���amG`����d7��!�)��v]�䈡����j|�v�	���rAB��#�Ў��j�cU*�";��l���C�ܞs�
�N�������*��ǒ���K��/=����_�k/l>�st}�_�8��C��i�+ 6`�� $��l7���2��͘O������QX;�_�+�`_p�hTU��ګ��~Ro�x70ś4i��
0A��ٷ��N�Q�&-av�v����(u�'d�Fu x%�u��
�����$�J��l�&3Z�z��hJ������)�e�o�(K۪���`;Zӈquh�K�"���7�)�#Ƿ��o�~�����u�ws|���λ��q������uL�t�#�`tKz��;�Z�R
]�8���Hn�>�\�9�j=$!5�<͏oY�3vr���s���r��FM������>Ն2:吻=�T��}ǞO��GZug��y"��V�Xr�]��3f��t|��w�)Κh݆��yE�c��F�Mm�^i?]k-��rT�,G����!�G��}��l���#<�.D'���K ��Ԁ/�����~p�|v_J�Yp᾽)��+��v�u9�=q*��J`EEz_	Qf-�֌!v���ێ�g�<uY3��^� �V�9Y�.���|��f^]�_e�\��6GV�n������\����u��yuTk瑨k�\���ɬ�mIM�m_��Z�ЗAw�x�ή��s-f�>`Ǳ���z-�$�f~�������'�w�Dsvg��5ۼ���R�H�J!v� =B	t�/�V��Ab��l>�Ű҈Q������|{���l���/:�8D|!<5jh}��:�)�{���f����{����1ҟIݧZO/�(���r2 ��#ȗ����L]��s&�R]~��i<G�'1����(R��LԲ�ͧ^���A��&풏!X�%�}��s�'�\�dB=�K����QQ^ ŐB^�U�����p����|}��κ������ݱD;ċ9m!�����o
̀.�iRXH�r9}�&���{�F� c�ݐ)��Z{�v��0�$����Y���d^�Ǒ��
ѻH�<A����s7T&�e}�0t� ��Ǟ��sL(�ٻ�e>Q4T���35G��qV���i��Vd�]Qsi-Q*p
��7��u;���ٖӲ<2د6/�a��"��/[#��zu���i������B�����`C�]e����EH�����V9z�H���1��#�.Yi��M���'������;^kvS�-�^��=��sBu*���#�#t`����Ɛl9Wŉ�c�����]��	�}W��f������P�%8
nN����m>���Y�����%7��Zp��� �BV��uj�MB�ĥf�Q<c��9�_�����{tqD�{6<��.6���Mf�Й�o�����Έ��G$�a�����Fcf��t����b���M�T[=Oib���Ȥ��Kh3�"Β��k+gO�އ{N�3��6�^�+�����/��&��>N3=�&:��;���hfk�dձ�D��G��X�����6�2�݉�Z��3�o(,�_�݋����E�E���N��1HUj�4{_�DT�`i���׻�>	D�58�kL�W��W�l'�������R��C2!()T�_䃜28R���(�h�H��E�`5��~s]��w��l���jX y�!u؃Q�)N�x��Z��Ě��o��l�LG��72�D��:�T���xU�2'���v�8�zt{i42�"�u��ޖ�.�$�c�Ŏ0��.��%օ��x�`֍0)�:��uT���߹��h�ŭ}�
n����, @��O`ZZ��d?�Gl�+¦�AU�i�t����JSX���]+��f��$W����>���\��Cݼ�u����ڦ�_�/���H�Q���?����F��R�`�2���I/��h�3+��2�s�L�\�`�;��S]q��=g	la�f��T}��^��q��̮k�����|/}y/TF���X�7�n{�5��wS٘Ts�%VQW��@��t�[�7�[�攙�#�Y��^Lt��6k��W@�NZ�o �sn��
	�f�*�'�iWO$�^���|��o5��E�:!�Q����o�VTV�J:�2�=����i�F��dN��������p�;�u�w�D��#�>=w�l^�:����E؍�z�D��?�-:a������ɺ�6\�� �zO��|���ā�v�p�Z�&@��mo����a�:W�pf�.��U��Z�P�лJm�s?ݰ�RK�J�`$0�� I#`q�6���4�HL�P�ض��$��fKh�	F%j�4��}�DrY_��Zy��qX���4e�é�R"�J[� N9Z2Ffg@��	�r��HH7�\��/d���t�����da��'����R���_vJ/ܵM�۷������[�x>���'�?4*�݁�z����	l�h��G	���m\3��sMq�}������ߪ֚�,�`D��c�E�gtb���O�Q��2<1�v$��@B�pu$-B#\��YL���<��|�.Se����X��A�MЀ�֕R���=�z�M��8¬Ԡ��%B@C�d<�ؙecS�E��U���M)�v"<��-��x�`1_�)H�{��ބ%��U����� F���ؕO��)^_kS�K�B2��ͩ���|��^��C4��R&�J�����R"
N�D��I�ħ(�z#��7���B�O��C�i������u1ݜ:�]�IcU
�jN1��nFi�/ʥ����|q�2A���e�����54��YF
H#n�v�t �����mg��~�kg��	�ɉ3��2��8;�caؾ[zn���yw���~��!��ȁ!�Y
ER�No*�+�,O;,�j�~�fL
[��6�5�������3����z��G�8*?a��Q ���I�^�ַ��T��	��\���>�! Q��.g�4�7��+@zrO6-�/���E��WW������FK��:���C�(���`���3	���0X
k�3l��<��Sk�m�O��)���2�0�|�<l�e9d@d#�4	�~7������A��^�|�[mPGz6�$��p���;��)(�Ȧ��&���x�A-�?$��<6�fݽ�@�<_ݾ�mV�)���'#�����>R�!�P�Ͼ�B��A�Db*b�W��݊^Og�}0���K/ ��V��>m�P����ƃ��VvLHn�ކ)(f�y�iG��L.Y�_��c�.�G5O��vW^+]��{�D���b+O�L{�(��� :�sk�C��lw�!��ظ���٭%��<z����12��4=���V;�4��H���-�.6��Re���U^#+�uR�?�q��H�5�D3d�B)B�<�[��CD�-L�T`+Gt�!^G��<�<���'�uMISO��K��ܩ��k�x� �&�%-m!���Ҧ��ޘ�%�J�v����nmyPR�Q�H���Z�~݂����L�C
�n�8��j���lf����� ��ruu� �P�q�&�W���c{K<����DDĸ�TP��5D�9�iCx�ɢӹx���#rb��&,W=�ѓ�K pp��ҝU��w�#�5��+6A��Ѵ2I��ѝ�vE�s(��?�G��P��hT���9w���|��A*����D!��J����#Yy��G�iE�niJ��YvmK���fܳ4QƼ�Yc�ǀD�RK�Y6�NGh|-�b���l�K��S�dV��oV���h%P��Q*Q,wL~Jj�6pf<q��j�)r�:͛<��'��$��I�0���d��!	�@-�-�*��^ E$���sN��w�≹��;O>��)>G�["�S��@v	�L�,N�Tx��9��DWokŢ��4x!ғ6,����g�!���.QL���O�n����� K�DJ}��Q�}��ll�㇅v�팼�ݯM�f��P����X�BT����dč0iIz�{l���CMtʩ�Wȁ�#��_3�7/v�پ8����]�H�(�C�D'�����~Pf��½E��muY�+/��1�xm,>�|�<�����ZS58�v��`m?�zZ~���J�nz�πCa)�	�At�(����?1[�U��5�؟>�%L�����d�L����l�)�JUe���UK�5�<� �>Ȥ�hu�KO���o���LI�ҷU���^\��M�� &k�j)E:���,2��4���&��!|�Т��Y�l
_��g�����I��3��3�:��O��9��Z=�D2��,�.)t܈�[�T���;쒾J��://��<���pWG�#p����G��xb�t�X�s�Z͹���L��F�&RS[��m�P=�X/��|�ؗ���� n���?��y4>;�2<j��*��p���?�^��GPH�c��4�9(�P+�k��x��(���q�����P�rԃB��y���;C{*���o	�.��35i+ u��o1��z���y�Ʌ�b7���$����%������?��`U𦤁j�1c�hzAt�� ���b�9q�#�����
��О���x���sUD��G�Oڈ>|�Z#��NW�FMmsA��� ;(�V��vf���n�o,b�gWQ0�託2n�5'7�@u��A�����u6��[�*UXXN���
Xk��R�z���}�����[��3�[�_F��VOh��,�'��� G�r<\��!�[ ��,�/ȭ0��=*�c0�ɏ�2
(���0ơ�C���䉳rδ��i�E�>�wx�X��,��c�Y�M Lo�h�~�/��u���4�fQ���+a]���EtJ��=���Ҙ	�`��b�@!3w�V���������&��?P@'c�e��K� ����Q!N��La5���:���Ԗ2����Dy�%��!�9�BM|�qVB���������h�sǩL�p�^ls�異L��S�R�xye��ԃ}V��H��8��\e Zَ1l���hytoӓ�w�H<��$��`,�.�BC��|�W��X�1T�qY%���Z�KE�>���ceR"|�V����R�A�ν�>�M%��Fbй��W�>D�B�q{l�;�n���7[���ɐ/	�z+���V��rm��[�#<��������Z:�Y�$��k<p�(�
ю�$۾��/(�^��	L'���L� ��TI���L�<5E ���n�pV���?�Wr?���×��-Zl\rv��M�jbK��V���WyE���҃ncrR	����\��Qc��.: ��&��*:����d��"��8af���oL\�s��ܬ�	,w��	
*޲�׊�0���)������5R-C}Yz�t��c.j@�k�������c�0�u ۓ��|q��?�H�;e��V~%�N�=M�z���w��.��k�0��r��lf�`;b+pXw����=]#�z���Ё�zq��7�'�`q|5�{#�� ����4:��e��F0�0�&}�.?�k44<�b���5͍k��^M'�ێ�a��%�'�^�Ǹ:wV�.���to�M�&p�(��O�n�
����%f�ⷪy�r�i���k^�_�I��0��@q$'b2Q��_����S��0{�Q/��i`[����#/�Q��=Iz��P�p� `Ck
�b^�C�ڂM$�5e_R^�_�c����B��s�?M>_�Z��Ztۻon�h+�[쮦Y��/�z�j�Y�������cT�@��ҕ�5��0�͏LE���mb�ޥsK*_���Z��8��hY�[��֔�QpE������ �r�]`Z��hZv�Τ|�5�t9j����׊�n������qn�4[M���Ր���>�X �ٱ�AA�:
>0�ŞlWb���(����@ ��l��d�.~�(�JЈ1`8�xW�Ȱ#�Т�>�ԷVF׼�t�_j{��1m�+��~e�I:L�����N=R����^>���s �!�v{�0�A
�42^@?Ń3���� �^#J�Sp_F1�6r6�\�X�`e���H��?ەP�����.�|l�GR�E�?P!Z1��*�U�Sc�A�D�N��[�����\�^��6���
����T��䓷�&��ld�s���[����z����C����+n�bַ�x+���:��;�������K�� W��qwK?�����D��g�^��7�V�78���`�&[vx5Two������
���W��9S�pe��0����9d��tJ������f��r��{%d�T1�n�ΐ#��/��K�g�예	Z�/\�I�����/�*��6��=X�^��qzg.F��;��ס�fvצ��fG���ƒ><3"��wW��>��h��F�j�u�I���� $� s@n���&6g�l�9&/="#е��JI*��̀nݣ��;`�ʆ��%���S:��W���&�_��W�	X��6��>��MsT�m޳ڞ������ӴB����34������5�$uD�!������I���<uQ�g���̼��}���@y�,*%:��G&=O;qO΅�U��6	�x:*���������D�"r��Pׄ���?�; P,�`����8�����l~�C]M��$�Ԟ�W`&H#�����bL~?�l���n<''��\8�/�3��EC�a�>2P��
��r�(�!��f�&[ݢ�C�2|�6���!)����" 몹�q�E�8�
�蹍
�U�(O�lI�B�B*<�Yw�h1w�&�f�tv,|-R���:?LSK6��}�dc�*K�&Z�߫�N���/��E�����Z��sY��`���;K���%~x�N"bs�n0�̚�cU/	ǽǬ�pvJk�078g{�ev���&c�d27�,zҰ@�Z
�㝎1�א�mg�c����Ug8k�:���h�
���v���c�4).?���H���q* ~���闖��P�bQk/R�?ae�1?�^2�������A��J*B��D�n����0�����f5#ppIa%4f��4p��D~~h-��yD��]�86J԰8Pu��8�R،���v�
���S�
�����ٿ�+�����\�i8{K0pƂAn�{�R�LUuf+������g�]��fL�G�>�� ��Y��`3����R�?A(���pr%JȺ����/� &��0&������| b�~4	bItg��A��s�i�4��Ik��3��Цr��8�R{	W��;jZ�[^�.���@9�n���{Ɍ-֡��57��q!���^�rY��ȯX��z�-31��ǚ6bx �` bL'�����Z4e@�����cS೸2)���g&��V�m�l��J���f	� b�ѕ�/D�;]j�s{���-
�p���/�M�*��\D�8��kf1Zm�z�4�`<��]�5�EK�ym	3d����v`���>�&��2��3f�p����P7����Qg 9���\���aj�Ӯf���Zj9I}6��x����O�+@rKA�TQ�,����
�A��wD]��>����&JHjg=��S�bК0w�(_��B�I�l��H���6dC�(�T��]�b��-��M��*XR ڗ�I��A򳜒��-�[̖:'b�rt�u����y�+�۠��Y�Ϟc�-U���5����9��A1�����k1ɂfg�:u�*�c�W����\�W�1W�>���>$��b`����^�%hϲφ_Qag�L��8�{SA�>��Q����q���+.��J�����WD�i�S�jh�މ�m7��\iF�Y��/#>�0zf��Q��0��q&�V�̛F�{�q�W���
�&��ճ
x���EX�&C��*8�s�*Z#�5͖���\2I��V�&A���͢���z����i(V�������$ם�g$7�^3V+n%�3d�OS�'C�'�gk�S��rQni&}$���M�r��瑊���_�+��M����n��7z3����Á��Bc}+�0�>�3N�]"����ۣrt'6�5$Bu��\jX�*�ٷ���N�[rlΙ��%�ծ�M;�f�{�q/S��Y�U5>L��;�lj�6�k{�'��n�I?�'p��n�q�5�*�4�ܙ���{fMZ��H��$��2�+1��&��/�G���*V{T˦GZt=��
��y�s�]�mo�ٓF-�|���"���}ke�L��Z}���r��v)�l����n�u����sv;22(�7�;�l�����&�#� ���(-~�����9�h�������K
#��[��SR� ��k.��� ]S���3�#��:��ܢN3<�'��J,��:*ͬU�j:�����{�0m��f��N������3
�y�;i��+GcLc}���'������g�!H�亩��k<�;���3��1Q:���N�ǝ!�*���Ϸ<���Q�eМ��!���>L6�f��I4
�sI��RM�����w�)�ℋed��C72(�5"M���{�\m���]kۖ2�"�tE�bT+�"JB�-e�5L$��)����B�n�Kt�����h�J��@�$㻐%�Bm�j�u�E��d/�� چ��!Ϙq��|n�_��}J��x�B.�Ph�s�,u����J4��LcYAyH���ٚ����?Ua�t��H�^%ߠ�N�e�ޠ�9��4�_�ՀQ/Zl^��Y��c�5x�`XlxVHYEB    5902     f20���W���0wҀe�s�K\�;�6�d����.^�{�U;��x!bA��ՠ��c��
q��]W
��tMY�D&�G`�{W!/� >i����믩�䙍�Ҏ�|�O$�^��̶��7�9�Z69DAA9�w�QI� �����Ӆ���Y�@�D �0�l�ճ�����DL�f<4	�s:7m�;u�5}ͲQ��'sM�l�)Խ�-��L�i�7��(���e��)�`=-�d7��PCnT��lȣ��·�x��Q�i�����?�F��i<tH7#���$�v[� 6|����� �m�y��eA����9E��ڬ7�2V���?�qY�!+��;Gn�E�z0��5���i<~0Ɨ�?Ǽ��U�Bǂ<M���sE1(mV�Lm�Cm[�6N�P#v�q6 8�).������"���-�{=ę��ze�4y�J~��J��'��>A� �|3u�<�O���iz�ɩ�K[�"c����8_�ё��|i ]-�U39R<�\��Rq�����bWKǝ#t�s���� �I����xj[0�Yd�c&Q�E��Q!��T`-��T�]+R�4�s�6�*�hz�v�/����t�K�ܖ;���cA��Y��s5/ݖ�tr��r�Y7ca��k������+�͉^�~��@aE�����2�����|h�/���=��Eܣ��
�4���Oi=�b���-�2)����\��[�	x�@��>g���8;�|���n�r��0~���V{�I^������
p�i�r36\���d�l{{#�6�Mo�?��ʴn�/���ÞR
$Ņ������qsVw�_�8�T�#�=�A�c����m�!pT�;s��r�+Y#��+9]�ۮe���n^ݍ�ִ!�gӋ�i���.a5������_x���l�'ak<�G��yY5�S��k���B�0����6� ��P7��X�h9n�o83�o�\?�n�X)z���+V��$���	{��y�q�`�<S+ ��ȗx�jr%��O��üNԫ����q�}��#���E���� u�X�ua_�v�mgb�(�lj��[�����g�s:C�}�6 �ᕀTܗ�9q5RirI-�y��X(wA�֖� �V̴r�x%o��]�*9�כ�w�ṁ+Q��aؾP��v"��	(����Mx�aZ^�g�@%��Q2�#NZ�Q/J0���9�إ�O�C���l;�fԳ���mf~�f���&ȝ(��o�ڴVV��>tP	�!�]�^�l�ݧ�V� $�`%�z𣶁�`������4�B"�FsE��A�i��~�����6��:���+u�0�F��	�8e�%��jn�������,� �7|_uX�x"j�ʌ�nQ�p�fiuѹ�3�.ċ2����Hΰ��LVg�E�脦��EJ��X �\#�h{F́�l�Lћ ;�^��˿�k��yE=��qWǳOx5��M���ۣWi;�i�Z���V���C�l�cW�rF�[��%E(xE�v�%�˾h&�"J�X�<n�a>d���y�$^U��9,���q�u���9���3����)��[�|&y���"��lߠm����׭e�e����iöZ��:D��<��M�B)p�?B
�Q4.���X��Ggyan�U����/
HEY[�:HbA�����t\o0�-(��2�p��9��S�"a������q�B'�������łJ]+��i�H��/b�^@�%�y���l|���!Ee��~�0�!�(Q���p��q�H���zU��jxvd��]�]'ۘ͗w��X���+���j Q�N�^��N�
RT q,K����H_C�uR��*�ĂԌ�8MB<�I(kq����r�Y~}��q�]v���������4�5�6�`V �b]�%N Z3m���~��wc���~Q~����uA�� d6��s�6<iG=������"��q��Ϫ.�GY��i�W�&ҡ���`��_�En�n(j�wKzJN�����g>SO�)��5�6-����I ^mU7�rT6���~�W��~��t�� ����X�Iآ;H��8܀:�t!��*v�=5�$n$A���z@��,��$�$�<^���	$���!n���ͣC �c��G^|\NF���$T�W/6�X���E�T�U*r��T��f�N*��p�2O�Vt�	B�4D�G��i7��R�z��BQ�͒p�aҽ�u.x�;�W�}9|��q�B�C,��S)���[�g��: �`���:��4w˚:���W�i
\|ݷ򎷧[+#�2�H�U��%��&]�� 0W%e��Q �րc��T����W�E�͎C�Xh�8� Qhh�P/?U���rPI������˙�=Km�'zٻ�&��\��J���l������)t���L�d2�7)(g��Œ���%E�j��G�ʽ;�i#��Wh�W�m���]�'���2��=�U6�xu�")L�}��G�d�"
4�,^)Ǿ��P��s�Hwp���h��כ��5q_��"���tn� Za�� �������R!J����Ωk��6��-�M���*��4��B��Zy�7��D��}��Vd������]�	]�"mx=�w�%T�>#�����d���9� 0dT]�2ަF�܎f�R�6�X��W��am�kZݖ�΢2)��[m�NG%��:���Yf &��fG����Y�������17�dh'��筨�]�$T��e�!���~���ޏ)���E����B�o�g&}g����L���1W_(a�g�΄u'�=}�.�����pB��5�q����g�v��C>V@Z�ł���J-/G�;�nZ���=��d�hQ�R���乘�'��"������,px�0�w��s� �OZ:=�}N�P�Ц�:���m83�&0G�%��D�{�i!%z|�eR�ٴ� (������x��_��]�u^���0V���j1͆�J��a&dH�뀉�@�O�p柌^~�+�!�[x�a�c�	�uIf���ED�BXY���P�����&�ԩ�/z�;Gz�G���������yȆ�B٣Z�t�~\3�X��z)���x�a�Ԙ��Yæ��11�D�'c�~\:z��sܑ�k�v��.X���.�v�@��4s�D�W�I�'�ԘE`#�T�R9��']����n�@�x�\��?����d���s�fp1��Jb�H���t�w��(+ݔ�J�^�I!)U��~�|��9(gL?���2����tk�� {=���AȲ��$	5NdA!}e	:w����l�V�;Z�^��m���Z�!T���q[f�����u'$`o�M��viN�cγ�/����7X�r��k�u��S���>�*Զ[~RӲA`["����rv8�<!����
���ʈ�7�}�+i���0Μc����6t--���)7i��^�o<[��� o�#ç����C--�F���L�V�W�\"|R�՞��&�1���Duq��z��ڹv'�`P�|��%����X-����#�j`$i?y��a��S�ϿV����q�毊o+�nY`��[r},�|%�dEw�Ï�*OY3B�G��܅�Y�0#ȫU�һ�.��ғ
��I��w\�^h�Ǝ�U�n���y�Z<n5����l:�w�w��rZ?=I�rt�����[?�H�-��_� �՚��O�W+�|`L��tN%Ocߜ_�m�N�a�M��м��u�oC<����+�Z���q�Z���p3
8�)�%����� q���Yg�_me �తeN���oZ%)Y؇��%9FcW0�@8��->�D��22��J�