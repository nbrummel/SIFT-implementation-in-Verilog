XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ԛmԝm�"c�Ĩ}� T^��ϣ߃��,�
.ţ��)�>��f]qo�h-����$Y���) M�lN.�F���oa!4�<�u8^����Ι|I=�V�ߣkxpu�4YD��R����z.����h�N��-������A��-��*�뛽vle���?�~�zV��3'�[�g�
p�s���a�\Cw�H&nu�	6�գ����Q��ߧ���P[7���Sқ��+�l�vt��a��@"���{�Ֆ9�0Q6���j���5y�6en���u�J��Ń4�2�ɱ�^۾�#�-~��*yΜǹgZ3$��N�
%ck#Zy�7^&��`���V��Y'�_��\�{�ծ	{��A�Q�Pը��(А�����Z�M7Ԕ}��q�iw|�X���=6l)�Ap�rɤ�),S��3H��.��,��sXT��7�;���-�ۻ)Qo��o5�T9�luPD���Rh���L��3>k%NJcÉo��=GgS.xO��ȁ������9��L�軫LX�Y�7�mr����ľ��m���żWt`�I���汭���նY� ��R�v��fm���6��<|�o���H�h>��l �����Hd~�t�,����EwlkoF�*f�XfY���0x��֔cM�H���]k�C5��%\�>*���EV�l=^N�ޘ��>�r�G�y�d3V��)���9���e����獺6~��ϔ��g�	��R��1�b
�=>K����Wu�+Pӻ�r�Ob;�N}I�Mj�d��}�B��vXlxVHYEB    fa00    2910v���dz4�u���Jxj>-X��[�ɋ�^���bT�t��E¿�^��SN0G��� ]~�w~��V�a_�'݀կ�Mc0��c���J��Sx/��n0�ք��|�y��~��&]�B����S���~㥛��c�%��9;G��dp�3^Z�^rl|�m�C� 	�+�X` �`�K�A�EB����M'��U(d���"�����z>\��{ T���l�����Ġ%g{h���L�{�E�u����1�q�<רv��eL�Wz�*�p����߀���[l)V4;/�q�LB�Wv�
���ے�A&=,}R\�Baf��纎��@�&�,�rVG�x�bÚZi�7�A��?��L�b`���4
ʈ�,�����l���_ �6_zqlh�4!��Ȍ�ޞ`Bbh:(��E4vr�|Y�.�7P�b==�uN\�*�͏#�j����h<D�_�N���3�&r�@	>��(�۲{Q�R5�=��F}����Je���Jn�xS� ��R��4����x&�2f��������AM.f䅛�H��˹�E� q1w��d���\U%�p�e���X��?��)�*�#S�6�u��D�^����lpD��._1�	�щ�Z��6���R�ilVr�����%�����莞�&5>O2(J�˄����U��a|3O��2e1�f�I�|���c$7��:�G\E(OO�;�o\�;�e(�E�+�*���%W!WV�[�����Q�wj9��ڷ�؊wf_������B*R�����7o�����j8�v"F��<_	���i��'R��Ы�3�����c��C�Ĺ��x�BOqyf��������X���	>�)�� ���B	?<��cP�V���>v_��`Hoh��!�j�)Çd����#�����f�;�@�J����i���ذE�Ώd�t�O�d<̈́��c����F�{���0���-����� khL�H�U���@Q%�����6(�����m�,Yf�4*��G�
�� a��+`��Z�7�xYW��-���*eO?��7m��&���(}�T#����	�u�Yrcg90��ݛb~�<�G(�I��9�6
�[�@���,==�_��A4$�e�D�#���Q(�M���e<YL,0wKe������7��8]���SC�0�^�5�t�w�I1wh]�S=?!�CҼi%���B�y�l�Nlx������o[�I���
�J��7cM�%��$,�bQ���1g��0��Lβ���H���71�~E���k4_�D;7�;��~h���t�pנ�G�������L�d8�d�m�ߍfW�A݁v�W).&&E}Nb���b�F�s`t/���+�_h�J*�:�^,��h�����;zi�#������/��x�j3�?8(���.� d�&�����4�Â��9�}l�{͞a\��uVlt��y��"��}��	$���eEH��RN'A玺���R$ɚ��:p�����_1�xD9ёK���`��r\F��~���C��g�k������]�3� ���E�:�9�]�i��G,���sI��hO�0YX,�U vioɚ_y�;]簮���ݯ����n�`���\�/�����T:��ԽpǳA	�Ž}�K�<߇�C(���8P0C~+9#�$�-�<Ͷ����)��+��y_��
��|9��mX�5�Y'���="J:==Ï��J��z��5�5�������8�������;��d�R�Zd�_��V6���������cZ�@����x���[��FA�k��>O��(8W1���ݚL���T �cc�ƞM#��Lb4.�f�����N;��d���?�����9Z��b�������{����F�zq�ى�Ih�d!p�4�����R��1��\G���.<�U:j��M �����|!1�!��_e���_����7/�RxX9f�כ����b��R=��-�&^`i@�Ϻc������NC9���P�9�8��Q���.=���\�����0��o��!�e��O}�q��t ��_�"��6�cX����U^ �����E*�	S��*�r�x��s?�{��m���_�Q����rd­c�I�"1��#�ϡ:�3�K;���gw\�6�d�W��OT[�����g�ڈ-LQ#:u��
�_2�I����̓�*�q���n_?��,z���e��,'r�"�hU���)"?p>O�|1X�Bx���ؚa��2)[�{ � ��d�0bP����Qa��A��BY����f�΂�R�<���4��,����.��@�]��&F����b�~c�[�"w/�eob0�ӣ��{"�c�1�/��D��Xh<x�	y�X�Y�f�{K�9ڐ��"<{�~��W�\Mq�Y�ѱ����9��4h�G�G�����N�l��G>��]Z�4,V�`,�$	+���ޛ�o�.�gyw��>`�pO:�|�Z¬�H�i�Й/���L3���V^ ��KJ���aO�A�)(��&���rSR��)==�P���zfR��������o��1>R��;�A냵��kQ��������A��-�C�����@u���T�!�&������oΑ�^K8�&�%UR?����F��0S��e���ߝ���Gk*�m@��LP/r�ۚ�E�@^�]�L�N�����(�� p���i*p�Ydp?}5�׆̰���K�	6���-i{ri|�S�W�V@(����YJ`�}5C
��z^�����`)���zM�-�+ʯ���t�ڋ�8��sN��J\���g_��(V���R#C܉��vk��E�� i��OU�~e��=�.���:H.��I�K.Ь��������A��*��P.�����	c����v��JTZ�JI�k2��ō��F�$q�H�E�EQ�� ���P���-�Q!�XL���k�U��Q��+یU�8��%�x�$�����>/�+m���$��]�U���iZ��j���2���t�g�;��,C���~_�{j��_�����#�y�ǖ�F��>o�В$]�
�jܟC����*��I���T&l��}J*R�Al�e�{�%�ѰOn�q��f����������zѬ1��\�_�T8��.]?�H����08{�0�9'%��8�S��V���]@Q`4�!}�iަ�+�-2�߸G�4j(,R��u!�ݼ��巊!�d�
��8����ο�뒷d�r]��:��ߓ
��e�Z���5�2z��bx�]�JHϨ&����@��q9�H �fQPx��}c�����n����/x�>W�囸�E?�mp�9�@]D�s��郚��3�TO}�ݽ9�P7��w�|u ��3�eԶ��o�TN��Oj��m~K���(2��ΙF��iRL�kJ4�Ē��E�A/skLS��ETbf!z�̬<[F��[��vR�]��]F~.��7]ʈ�5������\�
��l�p"X�q�|7h%�AS(�D<J/�H��H��{8�zf1��6 K1]�y��M��8*q��7�sN�U�!�k�Y~L��s�v���̚".U�S�I�(�ԕ�^/����
�Es�׊}Iefi_L�?���l,��c9��@��CE����3,΃_�EgM z���=�M�.�x��yOg_�5f���+�SmP��� �X`���;F*2��E���&���L`F{Q߂G�c>��@4W	��	F.�����$elS^\�_>8K��I���dO�c�qp��~����1��T�>��/pKE�=9&��G�bW a�a��Z�=�c��6?
� -�s�xE�n��j��n�b�*������3�ΕF���̴�*������簁�~��Un�=oa�{sTE��L�}�f�.
��~>'�i�
�Π�-F��6n���=ͩ�I��并_�B�g0u��Ǥ-1i$��cPa����yj�Ê��:��
'}�;����u;P|�t��5�ެ��]7�$��Wr�L�]8`���W�N@qI�Gf�H���:x
ݳg%{�D���a��|�6����sN��@1�3},'�a���P�4k�E�4��� �i
�@(T�����`�?� �
�;�H*A�B��w���F�N�������W��k]�,�J�f�o��}|�"��~�I��L��1<�BZ%��3���igQ!�f�a�߹�����d��I_f��4����~�H����L�f���)e�����k~�׻7���ݾ<1#��`о@�=�(* ��>���m6�`����z�oL�ہ'Z�������R�iK+���p�$�CxQ�첟d;{�V�� SB{?���d�X�hw67�>.���}O�Θ� �
a�ٸ�R�*{��jV'vA��K��SIri�}K�N%zΖ&2�>�'����2/�0�XX��\�u��
�yiϗ� ^>�JA�`�>����<p�Jm�����f+�MJ�'�j��2����uז_jR��.ߠ�=��֋`�5[*
�]Fq����� �=RW��p$�ilڋ3;�|<�|�G��ʫF ����W� W�$��ǶBQ=�Zy��T���Z[en� z�����|�(�T���@Vv͊�V?�/H�rH�	L�3<��zc��� �f�N�e���+f\w�9`IQA�A`O<�bڈ5&SY��<e=?U�mss+��<"s�N{�,�03X������y�ѫ��'���	];�)ѩY��︢�É����M��s���_V��ᐣ�QR>��i�O�%W�@"��67�=PJ_$�-���M4.��M��<+ �q5���	�}4U���_�"�ʓ�0�w�TkC��^.��^�[�/��˃�,(0A���nݗ�G���1m��=����n�3^tT��������D�l��;H\h4��ؘ�0��n~���f��JU������~�"PK�)lF.�C�Q4��F?�������8tP��E�Rb+����H�XG�:YO.Y��Zփ�^i�|��U����\�21�j�vqx����7YK�V���(�^��@
����^@+`נ�~aJ�3�"|��[�Vjҡ�Ȋp2��s��,������qW�S��j�X��O�B��������_�R�5�ce!`�$�%w�w�n]ծ�`V�t�jZ*�<�ߌm�ªA&�#H�.�3�m���T��l�R�8�����fqg�=� ���N��4�A��G���˵H�v��'%SЁ�yq�e�HB"� ����B��O	�������)@@�>B�m�eqͱ�R�F�[6A�[���Z��/B�txrŵ!�1-'4%�i����	����L�d�J���@�2�L%rJ�}� �Nng�9�=��$�����Ұ��)�D<���=����bE��~��E!�+�Q,�v��x�UWR��]�ށ}��t\^�-����u����^:#�x�Z'��+�((=u�v�av{�P�+,L+\E*"!(h,nj�)_���>c�h�(6��{�N�	@��}�rP��X�@�<G�M!��+��8m�*7��R_�ʕ2�"��#�^��#�M���
�
 �A�y�RƕqR�w���!��?��F�ڤ��#C����j��޲DM}U�%9RA�g�n����|�,��n�W��ğ��D�A{e���5�Z�`#j;��Q�[	���ܭ�6��͈�'� ��Xj��띲���t�O{���߂�Υٕ�:��Z�(�m؊�6�r_w��L\/�!`L�U�`��j^Dč����$0�����b����ED�>�/����D��g^֬T��>��Q�)}mȋ���E{�c�g�z�"渰�*i�q�ǝ}X�/+���bw��A��MM�<e��@d�E��X�9+��'������h8bȇ2v�H\&\��.��Ѹ�QV� ���Φ>�`���|?��g�{i>2��p�e�k7N'����#>P2�۸�rWD��ŧ]����1��(�,��!'khm��\�0�|���U��~[������,]+�XX�w��3�C�_�po[ԾwL�g�D�U�S7	� s��4��piu2l<l�Q���8&�3��(�+�F�L�r���Z���1��±O�lC_��/�����J���YQ��d���(c����,����6QL�I�5&��<���D}{u�d��0��v�-H�P����d��t��+�Z�2�ި�d0x�	�A[��Im�s���[�����5}<�B�0�(*�	2|��9K��]�~�vy��Qg�7��D̿�[��_z��0y��ړ�4���je�\�Gڒ�93�W�z�� b��S����D܈�^����'sϟ�to̭�A�sNww��.#�ק���`����JQq{.��)*�]�җ�Ӗ��<@��~̛�I:�ly *�Y&ɤҫ�b�/H{4]]t�T�劘��A��J� �I���\^�s���L��D%p��Ǎ_�9��E����п��s�z7��On|o��g%f%G��[���E�y��~Xf2 �i���7�?_ݰia�$��%��.���x<3ѩ��\�vIb�9ƥ/�u�&�H��;�@t�.�C<��4�*&80IC&'�6�%dL����6���.A�`��C^�&��@-�.���4)��i��<��e�,%(�^h؉#�}��'`I��6t�$�:��ȷ�ux����G��J��%�9�,s�o��Km��^Ĵ��B��N�{�r����W�g����H��)b���)��o��>�3g����/��0���fE��*Ԉ��_�K����$
!/8�^Og�MF 64R���k��Pj�/�&���j��rz�%7�Xg���3�{�q�(Smw�Hzʴ�1`>��څ�U��Y�Z�f�40,���� �S�����Q��	R����o�	y�x��,����1���2<�G$N4����-B�I�L@��#(`E �����W�c*��'{h����
����q���z4��`�u�R�Eڅ����J�Ť�C������u��_SC�'��h��JrB��
�%}�n�aD��M��LNy"�iY[��&rphJk�A¬���-�ij~�m9$' �bRݷ�E��FU�����F�G忘��M�C��e�a�����G|D�%��x�b����ç�R�Z����_P�[���UU5�}_�Mj;���&&@K\��3D`*?0���Y?k��g���!	֪��8��uZ�i{K�bf<�\��-|!���˰'�����K���t�#w~�-�D:�� ��2o�5�8n�+8~�[�UH�4P��v��$s�8t<h����(�S;��'3?[n���&�ΎX?��q$��:�1#�4a��L�S��A���*�����2�G�+!Yu�I��:6��:���ѬT�rѾ���(���AGc�\�v�۸@��Lė�i����N6w��@0f b�n�,'a4���_�i��pl�`�����=���Rh���f�#�)D�ƪ��lT�*��^=i}�������������r3��kPdv*��%���o�V�jl`y�8�Lt$Y.��J�:��~�5�U���Q�MG'����`@�'i�l!�>�}�����T����Y��j�}�J9a�Gu:L�Gz���;g�%�*P�
�4�����`�ZQ�G��t@Q0%�a؄9Z�19�iP~�x�<�"
�r����@�i�����2>ƿWfʷ!��}O�\0��&.�#G1�x�qU/.�����0��hע����ik�^��Op>��L��Ҿ@2���\�hB��B���##����t;�%������\_���G��S��cʰav��c!��ڞ/mݛt��^�U@yw@�)�SO�1V�$�:�)<WN����N�e���V��[vv�0��=:��d��yTP�=��6�3��.���du�����^�eB���/By�P����,�a{�^�OITs?��-?w"Vs7��n}	3]�#9�G!6V���e��@��|i�X^��mK�/W������Ci.u���C�D�0���*��I�zD�E�};��B���Wz�]s��!P��Rݐ'6B�}���&&x.�@릊_���L�_s������qF	%B7��ч�����f{%f��iG��#�d�Ar`�Q�7^���D��݊,�.A��&��+!�U�u'��g�ӻ��	�
S�Qu��h����e�0l)�����G���X�sj^ˏ_��0N_N���A�gĨ-3�J����VQ�����lҾ��I�Wne~>�2]�n�*�/$��Kk��{��?iE�[����l��~;��mp��+I;�H�U?�-a�;a���-3�OrX�0�x�\@>h
ӛ��<GcSb�T���g>=&�z ��e^Y��s�p)
&�ڂ����r��-  �m�˅�{�1��_7��Ӻ���g��ezR�Ȓ��j39M�Ҋ�;������h�o��h��5%j�^�Υ�LCԮ�Ͻk�JBg��m/Z!7Xq�b!a/s����'�r;�>X���8��G�#'+�"����.��݅��=����0��zr@�vj��9�_hc��3݄
g�h����K��A�����';��M�;0l� ��3�a6`�@;�dr�9S.���0;��^���-����9�2��^���bzf`�.A�!�ib�B� ��<e�L��d���O��H��#����$����V�QK�v��YȒ Y�r��]�C���Ӽf���U�W:K�e U�K�<�,T�\U����di&���OFZz��Mt��̼P�~j������Jj����=��2��a���W�����[�񘊠�p���O�A��࿹h��0>T���t�@RC�KX	E`~?��s��������b�a���+?�10�1ܵ:4H�H�(�fa�K����2�Z�`��ܝȌ_n1��iؾZ�V�h�@�9*�Г0��v0|����:�P+&݊Oo��,���i"�ߗI֖��y̹��'�*��V�qˢ�d[٨�<g���s��,?%�nz���*�`*/����	Uf�ܻ�ꉁ\Wyij�JϺ�)������GV� 9�@�3������KO��1d���Q*v����(�6{�����$�]^��X_�Ǵ���$�+��4��<G��y���q#������&�Q��-�BO���Q)�rL�`/����xtc��<�I$���S���@f��͠Nv��`���x��	]5�L%���YNe��0��.0:�����d\�������o���FY��z���V�L�p�v,�׳�kIm.g	�����Tʠ�ӕc�naH#N�@�'��Bl�C�x��e,���,Z-���攕�3m�h!P/Մ�'b2�z�cX��;�4�f���bfpea���!?����B�_��%�s��r���QZ���^{{t��h���%@ܣ���^��AҔ0{-�a�I��dÔl�ǥL��c~�F�oÔC����.Z�+��ҼF��-�� ���d�b����[S���$v��"K���S���D\��� Ø޹��t
deQ#��7� ��$%�A��=o�%��9� 4�^�!1��``"V�A�/Y�qH�m�A��q��˧��S��F�!�-�� Lf��>���t��Z��H�{9$ B�"�X�VF����R���v�����G���x#=���b�c�y��9�(;y�>&����]�u������[֝9嚽w����ph�-��T����|b~��	�V���-;[M>�7UY~P��nۗ2b�{n��C�^T����{z��U�F��6���Ҷ*����_�L�����:�E�g���/]=��u��.̄��<���cXW��ЙF��!��lU&��h��f�s��"U>���fc����(�_�ݚޜ���w��ʲ�Զ�Z�q/�Tl�P""���H�d�;ھ�����Y����-���'��7E���9�p�+�v_�����=}\@�IK����HȋJ֙+�#6��0�G���� �-D�*Kr5�ϰ��6nL����l��7���,@N`y�>��`&�k'�{�0:�	9��J�<�X��L_5q2F�y��㩣�/<�?�;�-Z�+�x��zg#Ŷ��>�b�[��e�al_g����r]%*c�����z#(}RK�&�v���g]'��F>�Z��R����-�&�L�Sb��������R�o@���a�-���O�L�c
�z������9�r�F�XlxVHYEB    6184     f80'����zn�e�$y���%N�`�
�:��ޝi W�K�? �)jC=²B��0��ȼ[�����B`�=b���}/x �U�y2a��4�h�-�e)���(Yȟ��'=�vХHB���>2X�$k�4(��e�-`~�!��4�p0!�E�g�ep#�
T�L䪉���)�N�4���>�$�t|�RM=�B2z*�3j����V�q�� D`���ӱ�"�8�4�w�E�sH:�XrwyY��(�Ώ��O x}�ca���D�����%���X�<�B�kg�}��f��C���5��}��^�xdc�,��B��s�Wk��w0zr����k,�͈�� ��"��tǋ=zQ� �9�G���<���g}���aU%�7���[U$�!"���7l��s�����m���|-J�D��{v^�h���w��GO'�{K�44X�������6֢r����F�Т�X%��UB�g�k��c�4�p�^8֗����� X(���!���D�yO��F�Æc��?Y<�|��1�I�2�\��ȩ�PM����"���U�}+�����5�zٌ���.P�w��2/DSS �e�z\��+���J�#/Zp%����1�S���5X����D}K�tѾ3��3݋��+�!81��J�G\��XH�78N����"@��v�&<�K�*�˰��䙂<�`j;��b��\�����p�t�`F�Ou�W�ퟢDd{"��"���,���'}���,�w�ٷ��2N^�<Wo�S�p�t�C��đ��T� ������KD���M�ɂ#T�u��ҽ3���J��VQ�s;��4�\c'�pX�z���yBi5IQ꣦��oa�3�!���+��[�/�����8��F�����T�ҋ�����^�
�����/e�iyu��x�B��ߵ2'�ֱⷩE5��(�7eKj<S�V�uȢ��Xg�'v.s��C���yCSѳ4o�s��ݿ���Y�-�i��8�K,Z�ԏ ��+W8B��\��V=��o'�ndf[�Z��ʤ�)2�w�F��G�-v/���o� ��G����_�2N�VW]�~Wf�~2�+�>�<WYsY3j���v���)M��3����`���M��N�!u��V�7v��ٓ�gػ����m@`����T'N�O�����QP��IWy�Q�|��UR YG7�Y�%���)��
���t�4��S������o����ab���������G��J�6���G�uO�ߨ����#[w5�4��{x}��Wճ�Q`sq�4��Y4�*{�Ǹv�,�Kk�c#l�=�?1DS��]x��j��Xi��Ԯz��˰[�kF���G�h�����7���5��x�j�<d �hId�����(��|��D�v���+�d�[g�X�Z�՗�� �F{}z�����r��_pG��N���&�K�w\ ;��m�.��H�߳5׵oE��n��r�B�v�������U�bk�4��@�fF��\�G�ZU���SL�a�����d�^�#�oj��>Gk���ϻ.��![��j,q�Ţ�J�6�wg��,��j�kq��jP�d��w@����J��@��������8�����w��]P�MVٛ5Z������C�x�yݵ�e`}����ͳ$�z%6��@�W؂k��u���<���m�^!��1(�?b�W��9X(�I���\%I\�����:�Dq�Y6Dt.ً���U߰>u{D�����#c}����5��߄�"7��oKSJ8���~�G$�ip�"�l�x��?Yo�����l�H��FOZ���G�BK%d��cC����p�~b�~�+Qq�-��G_\��]@�g��A�5���M'K/�U��'��g,a�2zԈt7Tgb��1K�
���|R:�c��8Ք��h���
��5;-�+V���v�Ƶb��u��9BE�?*�d�ɲ���Q1{�f�L�#��J�}`���s·#ߙ��u���1����`�����Z���d!�y��Iw�䮕2�*
�q�l����D�Y�������:������y'��!�G����)��y��pD�j?8t�z�XC���%a���*��%i"+�
ГH{�e�>AS�/�c;ʿȊ��If�*����9����(���F�\��![��?ނ]��]c�������eU�����}5KJ���W��*�U�-�� ��e�hp$�8q���oml�:��l���������0�W�~& @�������s"�}"����E������ِw��/�hy��*'"���$ ན��W�E_�5�,��ӿ���x6��nj���2���_�(�a *�]�w"������x)e����������x�qk�;�\&Xƿ63_?��j��,��|��Lv�&�N�g��P��<�&)�1���V�kú04�c]��	��nZg�T�������ө�+�[�4�!>+��Z	�@h�
�u�2�h��-��Qg"k��(d�x���w���`ڞ�o!c犷?�CH��I�~=�^h�3�CN1����=QW�+Z`��D�E�yJn<�p��gQ�dmn�VcEt����+-1����6�G����R��\�"��Z}4/=sQ���{�2�Z�N�c��\�inpZ?�"���n=���K��b�j��Y�HR�k?Z�NL
��4�kU�]R�O�Mf�G�2z�:�o�f�^������ �6
�	���1�����L�����c."�U�.�N��\Mlk�9q+��-�8S�H���lD������j0�T�'tݠ#��s�]/cU������dZD��ԧ#7��0%�������G	���;b��U����o|�]96����r/:M�,�R���@�-H,�����R0�P�S����6t����?�ݪ�l�����Z�}��<M�7��M���2|��^e�ý�dA��熉>�
�k�7�u�t鷎̙3)�P��P��44)zP\�����E�B<�j�4�8(.J-������E��J�h�+�Ì�G1\$�g�	�H UD����eg��LF95��EN}����
� ���ן��[�9�O0g�qD� Z.�M\{���K��L�jP���I�@�&Z�Z+���cV�������Oo�M�زbA4���nEY�!��2�C�,C�ߝS�����O����Z^�\'�~��1�v�o�<����z�8*�������C4�.E���(@qD�]��T����G.��`�ƈ���N�B�����^'�:]�y������yC��Y�b��1P��O~gH�m�n�������V5��h��K��vܟ�Y4Xj��~~"�V����d]{gS�����^��Ȟ�t�*�Qq�e�Vb@���y��Xr 㑉a��V�ǥR�K�2��hq�@a�t]�~c�(8
)P�X򕼒>�V���tIA#ES)�(4�[�]��L�w�,��z��Iv�D޷�3�z#�Gi�����0�7�Q�e&�n�y�������
y@Ʀ*��E����;X��7�
Ԙ%r�O�|��Z� ���}�fLA`M�у��^I{t.�Q�$�7�>��dT�8���TYk�\-��Hr��	�a)�/pAf���w8����ݾ'h��[�v|���o&����ê�UD���u;kV����
����b���**�X�{����v*f�ʏZq�#>U�*��-�k0@c률�M�>|6pj)���W`���"���
|�ġ~a�͜��t�\Ɉ/G�R�J��t:o���Dd/vz%�tc��|��Y��-�:s�b����Z�t���,
pC}h��%H�ڴ���HR^k1����s�"���3���v�����H�|�	�,)�2��13�[D|���R�z��g)�B��.�~��6��1ߎ-�_82��h���[��