XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���)<1���baj.|S��!�1�'�e�~�F	��$A���.�,G�{����rhĬ���g�ܜ�-WY��X��EqȽ)�pm�	0իFtL�V�bL�����\�?�l�DA�=a-6�d�%��Dt��4�QIm9'&9o��ב�G-H�&����Ƙ���RU���9��՘h��E�u�B���%�`�-�˴��}jM���Gr��bi�f�T�������?zɂ�W���]�_��d��7 ��Scܘk�r=�R�������R�Z��ڔ�·r�gycTH}�Rvt2�P��$�@�i'���`�C�yT5�o?��w�Nh�o�\�����.��"J�Ř�L���(�JY���xeފ��A�w}��ɯ=߾ྦྷ��U��P�M&�ވcs�
N�4d⼊!v�|�!�\�O��&������<��� lƛ	Ktʭ���	O�Ч���1���� Ci"V�Ky��.s�D�^��U��4<K��Q�\f��;�.����A�h��J�Ov���h�2�-K�@u������`�����˼�g N�?�;X@9bR�EM�C�ܨ���3�%��6�����g�	+�\�v��$-?X�A�R�p(��hw?�ꮸE?�-=���l�آfi���C����X���k����Q���_��S<��r�\�!8��\�0n.��wl�J��#r6I� ����7L��.l���a�뀥q�HM=ϳU�|��W��6���XlxVHYEB    37dc     af0j��i�x�a�F�z�9�	�A���M#��x���
M�!~�� ��4ic���=�bbc����ꦠ�{g�*pI(�
B�-x}���y�{l��߷:�PeX�Qf���ת���G&�Q{��x]��%nb�rnlm�7���(h�H�x�*�OQ�Z�Qv�]+�~����;�>�<sWB�,uo���C{�6�AH5���H-4~&�D���tԏ�5����*� �<i�k��{j9Ԝ+��rkW)�V�KP� �9��zV�4�ڭRƝq4�Ǳ��V���
c�P���>��D�8F mZ�VϺ�Ǩ�=7�5:oԠ�h�xA#c���ϸ��#���[���i�[�����׽���$�I�J��o����S��x)x2b"3j� ���Ɠ�d��C侣k ^u��8n�ǭ�f����8���c�����,���|2�������Lc�"vH�j=T],P�Q�]��Y�q�Nv}xƨ+i!�=.6�6v_C��h��_e%y�-���o����x�Kpt�����yto��#7p��a�o=���Wv��S���I%\$����<ݕTYZ�� u�~[��rC@k(xp��]s�'ZO�\���x襦��$�K�,���"��j��O6}|��_��r� d;O4�~�Z�z�1}��IMS�ğ^��b�϶���/���eʃ�ip��H�MѨo�^E���:rA)�^Ӧ&��F2�Y2��[�b��C!S-|ec����*k|�_W-{j�ud&��bo�XW#�	��
0y��V*�!0^H#�}�j�u�����t�iA����s@q�MH{j��v?�����4^Eӛ�oW���G���R|�K�$�(��I-��^��_��ѯA������۳X~/��u�j��h�N��`}����e��,�� �x�����.�|��F�B˟�xI��X�ب������a���8���>9�Z�f+jt:=��e����r�[c����7J�aL�ʥ_� �_%���!7}ᣯ�����N ����PH;W�:]v���!�cJ���C�0	.�_\�=�##��6� �!]c���7n��Th��X!�@�ǡ�-�6^�IS��🃨aߤ܏���sq}~N��3tJj�6!��sCFm�LP:��:�n�4�l�o�K�_�Y.		o}�\"�"Bס�X�|-_�+p�j�:ʯ�9�f�2}|V_:�҄<�
�r���{�1{j�ڵ��_��ql�"�_��ς����Y�H���}O����P����Sb���fɹ��y�B#�t�EA:��)*��d�:=��7�!�`���@Yf�Awmz���J~�(h�[�����F�|��\#'|F���1!_67mJ)�|0;ЃE��Nb�V��%~�mʴ*��!�j�gaC��f%�]�������mNR��a�{��ȑR���޼�ft\V�g�Ө`˭i�4�`���`��5#X	N$f���YvpS�
���]�8�����E�S��(��:7������o�e���_.�!3O�ڝ/w�h�J�����/R�E�"x8�9�g�*pfM�ʤ�/S���zh�����tx{���2t�a^Nβ��U�Ho�D��cR�0|;�XD@t2�K�]/,)�B|���E|�d�p�44G%g�Y�~��V|޴��|��q���4a�����o�2@}��+d��� I.�MǮXq{��@ٝ,�H09@>�s������8�cl�*���ʿY#	7֕���^��n`�?6GOJ;����8,=@-�,�8�M֌ɇ�x��?����a����ӏŽ����Sy���Z ��rE\���M瓧`l�~�� '-�B�6C-V6�:�����=]���|id����!�{���4�4�O/(}��<JԆP�.�3�t�;ra��� fb�!Eף�i_�u��E'���ݷ'D�u�����c�Q�ȡ�}�g�h�9ɒ���c��'���B�H|~��u���0�:e�p�eg�OǘD�4�l�HuۇNQ�� �|���es!!�CH༳�[�����\R�2z���˿X
8x�1X:}�#d9m��W���E�M��G�^��ue��O�"Z7j��N�����gV�   ��F�ǘ�O/��pj�_faFR9o�����9Mԓ���+5�f�쒍�B��x9p	���h���1�4U�j,���6��,�V����#n��Еx�(�
و�H�A�z!8x�/��ؤ#��t	��up��_���'���Լ̪�����=���<~8-�f�ɧ?^!���5�Ӻ�١1g,N6ĳ�r2�t<�������Ԃȳ�S��o�=#�m�,< �R��n�Y���՜lZԸ;_�+]���2Ut�����)/@K/�	�$jz�����rcCT�g�-K��8�+����9��-��AOe65p>�Jna`~8���Fa����c�lb�Lv���3dF��ݍ_�qV��� �����HN"ٜ|������{��d"���Q�de�Kn�8�w�Ct��{_5AO;��ݝ����o�� �G�}��Il��@�%�>"b�t+r;gl�ş*
.K��Y/5�k�E�I�����{4������	�S�1��-�t�?��h���U%�'uI�0d�Eg����[�L�-��س�#������9O�˼ݶ��~�z�\-Hk���X��x�v:b��t&���A�]�����ص��RK�#oz�_�f8e�(b�E�6��Є�����+��L:�