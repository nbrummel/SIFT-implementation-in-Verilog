XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0�K�y�zq�z���8�����N�+g����̀�U��ڮC��]df����9(���}컧Z,�@��4x݁�X?Kj��.�u����g�Xh�}�%����y��g����Qk�4gIo��0X������J:���]'@�x(
�p3r+��['}��߈d�Ӕ��Ji��:�������X̂�Pt?�
�,b�����nl���JƂ����;ѧ�,U(k�J%���_q�_1���^���U
j��֍��/��!Sʎ�m�F�K�����렧�7n��3��;}�<��G��5�_O��2|#����2�b�x�p8���l� �q��ʥ���'��7�q,�lqrk��y�@�J p�FYI}x5s?<�#��wa�]����
����H�
y0��Ah��3U7u?���X���J�g�n�d���o�ѧQB�#��jD�3�cy��$w��xA�\Α����LCXcF~m��!�U�u"�B�w���<����5]|	��D�&ٶ��k@J�:�bC	�㳝I-KKɜ�5(ϔ\������6CR��)JUt��ͼ�1�!����~���Q�+����ϡ��{�S�m�95��E�X� ]=Bg���#�t�7Ð�^�
��z\m	��f�.����J��(;���ϙ���Z�y�U[㓫f��h�u�`���w�(�p��kY}�^~�?�>Ҥ=��c
M���"�.݅���I[���(�@����$�����7<���4?����ʹ2'4eXlxVHYEB    2a94     c70	�$�ù�"|P��[��^ZJa�N|OF1��*�����9��xW4�b��{����p�VUV-����HOq��C��2�R����ROŇ\�p?J�[�7�h^.8�U!��Oܛ�l��n�C�7T,@6�@�������b{��eϴ� ʰJe�	H�Z�Ju�#�|̟aNͩy��7�3J>(D�_~K��g�C���{���Tw?��=�~��b���B�)!译��S\®i��EÌV�X�����������\�)�d�e^gT�#��#�l�&+'I�	xw���}S0�N@5�e?T�Y9����� �}K6Ϋ�sZ��%��I���_��m�%U0�b�"�F��~vL�wO�{�����$)�%���p���A��I]�-<G���`��d��.��r�j��C��2`��;��@O�_+����S��*	�7~��>�E:/�qU�I�%2#3�/�q���^0(ʶ�T� ^aTp�jM��#Ҭ���4�+/�[H�O|˙�Ma>�L���
=��=��* 9�e����@����`/�3��c+�4ߥlۨ����l;�M1��yJ{O�!��-�#L���*�G�8S�8�p�έ���q@Ixd�$�ϔ�X�I���@3)T�/��}}|>_��9Y]��� S��ɭl��{&R���bV���
�d}�>J������k̦��G�p�� �M]�e5
Huq�����b������S/��h�{XB'q�o���S��5���gYG�g3rTvN�{�&DT���u��1���nk�hL�;m��D�s���%u[	R���[�_=<&��~d�:��_s�kRG��7�dA�I�uNK����Փ�qȯ�����{T��tm�?��in2��6Mw1�K�q�3o��|�4`�F'ҏ�;�H��Yl�kV���q
��}��-�
`��x�����8�F�����( �<$��h"������o�$�n�{�7�7���v'����@,�F-f��Q������/ָ)�4w���@��bta�D��v�Āv����k߷�gmKrЛ2��ƙѢq[����v��!��[֟�ɝ�fDk��>7Z��&�W���}`�o��l����ڹ��Ε���aj��S�2֡oQHV51u$C�
>U��\��bz���)P��d�S���z<��c亨���FW�9@�oFRֆ�	��T�EEЬ��_0�
`�3�����i��@,Q��;���B�oz<$\ӛG˨DD	���To�į$t�^�:����(Պ���TG�_�srj�p�Q�2y�x)�Ov:�~$���,�*�:F��3z�~&�S榒h`F1�f �e����N�Y��W�ծ�~�=v��$v2�v�����+�sDF\��~1[�K�XȁLӤoH�\�=�� �T����f5�����B!��B9�5
x�U��Y��*�f��������s�l8�+˟Q*�:G����������qL.ȸa��K�������OxpC����toI�Ae8o�#�J�I}��k������f��J�fK�AFZV%��D'��ro
�i�_ETK>83$J+Lu���N=�k/m�s��`��!(�[%�˺�B̰�h�$`'�Gn��`���	&����1�2'ί�[V����\b�K6f�����l̐�NJDI���F�S_�$��x�~�;�޶�B��-�/��͞	zȤd3,�� �U�Iz�p,_�<�=��ݘ%8�1*�������Z�Y7��VW.��c^���㱑�H��]��/R~�φDn<��M�5���[��c '�>9�J��B���) u#�=n^���R@�T.��;�Yb���l��9�Q��~��r[��G}�t�0%K�G�Ȯ)�c2�g!tm�%�����[M�y��7��{G��*��C��P9�4����u9�.���"��7|L�Ȕ�4,E��x��	��]%�S�,�y3!'���6 !�8T8�|��~�*����a����������b&�/�H�O�69���"n�}���,Z��3��t��l>l+8ChF��3�KU�8Vd$�AX϶��}��|��4M*�-E��,�LhNe����>(;.�g%��tg7	��̽�IH�Z��h�a�T����%�������*�5�z�X� 6������Ee.�{�m�&���s����T�:$C�<G&u�l���,!������+���w����]�o#-�"�٬0wVV�OĒ9��Ϥf?���j��_�"�͡{��s�w';�`���O�8�3!VM�0��[�O�-bv�Oap���1KҴ3������M�\-��9� AWw �YK����CU�%?7='F)�i +V4bA��kwG�� j��?o���	D��{�ӈrQ����>�_�F�����)i7u$��k�j�J;<����*��@��! �����p��@)�D[�h�p��ȇ��[�4��<E���e�
A����k����XWR;|K�:"�/�,�O�='ZHk�����+ǜ�N�|bh�1	 ���e���8ʫ�x1Iaw�j�s�Ԓ:�n �FB\,�{6ѱd-�K.5����+kl��szsG�}�)�w��[6t�+;���~=���Z�\���{����\	tWjbdQ�Jɩ���áx�����"���^�.��� ���U�u�ǽ�7A���C���w���a!z�ǋ�z~��7�BsWjS�~��v��PS ��U��Q��`�R0�QQr�'���jy˺�;Rk��6���;�����H���Kj�����!��� N��Y��!�=��?�D�n&O����JE�*�]�j�k���a�f�0��bx�-,%�4+�ʬ^�SPZ#v�u!��>̙����檫f�`����i�G�C��Ǣ�F,KՆ�V��ҳ4��yT>y�lW���T�7 QH	���@�Lr�`-�^剨���d�������J�fF�s�W:���������հZ-=�XZ_�t��7n��Q=�cv0a��_�9AٓSh�e��X�`�g/���=5�i�`�7�������b�X˙�,HK)�(g]f��~���B��_kH�Yp�$F�����5C�����a��qD�����P�)~�o������~V+���ՙ%���#��/�9x��;`�ѡP