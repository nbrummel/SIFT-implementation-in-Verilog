XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���24e<�ǆ����yA�;؝Ȃ��{�0Pk\��������͙��T�g��b�"��&Փ5o��>T�^�i7Ґ���j�f��]��[J�����w�l��laƹ\,9�W9��q�O�L}fC������f����R����ƽd��3���Q�^N�ם�0�,���L1͹ĝ�TU���J�#����l����pB>P���$����E�4G��iA��=K�_�������}?���sk?J�*���F�g̷Ȝ�p�B]��*��m�	�2#2�LJ���t�j$�����.7H��V�@��D]��JΡq�oķ���!�Ԫ,΂�D�!�c�kc�q�ď�I ; �����]�Fs�Ḣ<�FjbnʜǓ��qw�$=�m���M]ъ�w/i�I"[D��|SѳO����@+��U�؇lGXb�xf:��+��L�M�*ea�B�w�Vt�d��C5:�H͢;�)�S�V��ѿ����;�?�O��]?�V	��o;S����8^X1X?�1�������*=A%�K[>��Vl(|P�D`<]^1X��I k�>�~;yԴ0,�ؐ��Lb�Ou$�	���F���6ˈ�WOԸ�"5�����YvR��!������n�8��&�_[X.Ƌ4,�S�x�+�a@��b1�Py�b��*0E�����P���Q���K�,��/	Sÿ��ڡV� �����9�?�>U�cP��"F���C��+�HԪw�n{���RN���XlxVHYEB    2dc6     ae02���L��&H��}Y���6k����UVer�"�i*^���D���2� :Xqd����A�y��O�fL���l��э������w�ai~9������h$&��x�����!�-��9F��[6qA��3� �`�����4�7����7Mf�p�:,BL�tQŐo�Ux9�c���.�������gV��0U��� �~F�
uf�s�~N���J�t��jq}�#��|\��.F��� Pqi��x#��2e1�ǧ��/Ǡq�.	j���&j��B��::51ޠ�T�3�u�	�7�,������&�c����`�vbX����y�`����Z�;��d�H��
࿭�G���-G�NG��Z��R��q:�R�p��/i��{96��fXT�R�8�R���ۘ;w��?YA̎��8|�:�uPK3�	S�F p���k����O���D��z�/6Fޢi�Lf>�AEH���#�R앖�ā����G,�ݢ�x�ED	�Ir�����nf>�\Im��夘x9��hP���'YQ���hh,)�eEc�G��0��V�@�C��9Hri+/�v�RT�^Cf_7A혲�qO���e��/)��'R�e�0�2e����G�:���%�N����;UEDֳ���twơ���`�����t6�I�h����#
��+���J�%3�i���ȿ2A^��������]�U�7F�>��@��~�M�.�ᰋ:�Ԁ��Rȣ���t�	��l2�`Rk�=x����_M���9X�H�jQ��p|{l��xCI-��$k�g�R!�J��p��Qh=�W�;��CWK�!�!�j�W���h.���ۖŖ�tq�sӦ�����x������zs��XO������
��%��j�yf���Z��rb���7�	���I>��q��5��'V�2&����!V�pC���Z8[8����� q�:_Un<���i>���oB��U��"��@�ImU�(mZ��X��ۭ9��b�ޘ���Q�p "i�$��*���-�gJ,���m�g�2$��f~��nH9#1Ex/�b���?!ܤ/P<�	#m���Q��\;9p���J�`6��C�WG��r����@y����W�c%���L֎�u��2�+E<��=a�
��1)k���֖�C��u�(0����x�;J�����ޢC�ź6�&Pjv�^x�,���PK�ƃ-�֡��� �J�>�Efs����=+Q�ؼ.g*&2�o��P�M���u��R�����R�\�>ia0]�>��y<�v�~ K�8�jz�� ��Z��;F�3�{���*꨹j|iC�/�5@}qB��A� �g��jB+S���?Ē�l�^������/L�PTl���Y2��æ��������oSt�H]��'	
�@"\�x٪�4k�+R�LD�](�ԙ5e�8��>*UF1���
�.�k�z�z(����2����x���x	㒭f*���{���`��b���Ԭh����=���T�]���t)?oB�t�<~�9��o�l^?�"	���yLꮺ:(u�N=P����coˤ�sT1>���¹���1����*&K�d����[g@�Ν�<�	^=d*�b����b�酢D�}���άqbo�$�����p�fe�wv��"Y��\�);�c��[��V_6�J�n�CM`]�J�2�e��4ƨ-/ۓ3.�.���B�b��Q��aR��+Ȝi�ٞ G��H�8�q��}$t�'�{�����!΁�:���Y�k� 	D�����a5�� ����k ���[���ϻ�@�v�� Y�~�5�k�`e�	��Z��s�ے؎���,^�a�.��&��,����']A%�L�������s�p�4�'���D�D�`#jÞ�r�f$�z���:KzĨV��q���"�>�e��4c|���3H��Z2��1U��;~$Gu�b�Z2�@�e)_WW���m��T4O���'n�KjL7���Z7�r���R�O%�ANk?8J�?~���)y�q��,��Cr�1�|ف�bp��J�-F�Is`'�M��~J!& �i��ۺ�%�]6���RPwvZ��u�%�򬺾ȗ�I$�/˭/�ma����[����c.@�<�����A���X��g��^�>�W�D3{F�f�D>����]@�5]q0���b�m���q$������_���2"�Mj��K��!�OKb?���!�����L+~;�#����u)����7~R�a��EXܴ����]��ߞj�
�5�?���<��&0�uX�֐�R@?��zǃf��%&��w��dQd_1�Yf m�9l��FH6�lާ����C�|��1���c�� �W��(k�2�L�E����E��CF;����x�zO���Ck����!0������d��OqS̉l�F}=��ew��1cpͅ{>�>����!�x,���(�:tq��k2�F�|9��
^��:�����e;���\>?z��|�(�E�zt�y8r��l���������7aV�t�%�ř �rm֖y�΄X#�uV |��bz#��!�����f�L�d�T 4S�f�p�ȇ>{U���Q��a�}�
2�NC��,@q4.�6�D 03,��@�ˍ���Y�WF�9�'�t�1b�?�L\O{b	��5�W����F�	���+�����7�5��܊<���.�Nd#���