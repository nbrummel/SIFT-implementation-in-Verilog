XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��O�
���i�t��%����,�7��f~�[�@-�8E.���*>օ�V��g��Z뿶�s��_���c����A:����l�B�b3\���D���x��x��K�~�hA�=j���	�7W�z�_P]0����|D����=�xB��GIb�0���&�g�mv��`��ѾD�h�I�!�-�%>.Dq����DێPY����Cn�o:��烗�ޓ�W���eW��-��J�v� J�����K�(4E��)�����ȴHn@��r�@Ow:�#�5�E-�_��W�6OL���U(m�F�zˊ���~���L�#��mzB�E/���N�9����P]5���:|�S��)�LO=����pj>��w\���՞�ԝ�jL���+��4�祴�U1¢���c�f�`i{����o�DW�r��<ܤ��0���A���[��^�ˬ�v�ݲ�-�b >d+9g�D�K.�� ��E*/�n�'"}�i�*$�Yuj�=4C��+�Ke�-m�6�o�{�y̍�8"��b� �&�І6e�؀
jӖ:�Rx.r�+Ôt��޶�r�����y�5_iG��
�u����<��S;�����3$G�,&�a�����僃1K�x�r������N�}�Xi(�{�ʱv�\���:�K��S SO�C�ߏ�)�ð_	�矛�b �T�1���P�k�.�N4 9d$5k��?e|R��6Ң�Q���w�|?��8��~P~,2[Cn�拺
VE�XlxVHYEB    91c6    13c0)gz"��֌1||����ʞ8��V*��o���;@�V1� 9��&~���"����&@����݃�5����G����X@��	4������
$�<���`$X�×��r��5,1C{�	�1���M��u�J�pF����c�b�)sx�j�akM�G�m`�F�ZT���Rd���5;�8'U�����s���t&O�KYKw�T66D���6�VY(��\�r0p��#�����*�Pe?��&ײu�j�3�����U��]��Q�� [����=U�i0Ǖ���N���X%�`w�,,�*89i��NQMpX*��Ah��8*�p��L1������H'is�ց�V%�%*O	��}ܒ�[�Uզ�ƪc���=�UT/�1�$�ƽ�<5?�ΊP3?7��'�c�����(�Y+���;�t��;o�H����7z�˷&�_���L72��'�(1������+��W�w��s�HM\?���j�Aݗk����!���a�s��ѥ �gpL��)�G�V ¶�Ruh���W9#�j�1N*�*��IDZr�N���P�����y�Ej���Ml��;���w^X�(��M���ƽ���"�ӯn��9ĝ^B���G!���r6F[�g4b��lS��g��:�!S�2��wb�y�p@Î�P�*������`rI �fwȃX<���I��"�>��M���1+��km���z�������|pI�C�"�lp����j-m�"��v��]�\S�T��G!(�|������\!/w�AZC�#6MV-�w0��l�SO��|�^d0�V���D6K�f�n+:�K�J �9�( �me"��8Z�����d/=�2�1I���+�K��ə�G��~J�����d���V����cς��	 ��5�H���wOs��.Ⱥf�~�CJ���:������=�Ą�~� ;���+0�tL%_G�=����[F��r�T?�����f�N�n$e�7�U4�>�����:���n� PP0����<S�O���`�(E���@u��& 	O��^摂�.6��Oڷ�<�`z3v��#EEǽ/F"{^����u�j��_����ن�q���q6�
Z`+�s����%K?��R�m�Io]+.��:�G�N�mYȜ;�U�&�_�m��~����bL
��w�����y؄	�����n�N��[����ɡ���=,{F3�o;!���Q��~�����$I31� e��scy9�"�����yo���2
�:\"I)+D.�b���G �pW���`H1�#$̬��q���)S��"�h��N���~ؔ��/#��H<F'�}JB���8��T�Z)��_j��������{K2���xp7_������1oL��!*�� ���l}Lbi9Ў�ul<�ya�z/?	j�#���'��[��#;�ۿ��LH��F~zȋ*9�������a�z=�_�tV`�``|�^��c�
5��Q�L��p����|��Pk����悼ݻ���F�m;���tt^��(�#{�%�x������L�����tʉ�h�ųl�y�eMW#;���H�vWP:�~�^�לMX<)���o�']A_'�k�V3��(�\�I���-g2q~�Xe�1������tt�YP�$|��m��G�ѽ�����׵����'��=�V�tߨ\08>Y� ؟B����������a郒"����c󹁙���ם��w�h��'�dF�)]d���|�F�e5J��Y?�">�^����w�1T`m4�ٳ�Tu`�v�y�)��.��)a����a�"!�S"@�� �y�X\t����m�3A��2n[�p�U��%�
b�Μ��<��@�.,�Q3��'����e]�<���'�l"��fB��q�o�=������%gU�L��vv��d��u~m���ҕl*�/�HR�y�F�Xm^�bT�B���T��L�����
�}��&�,�ǈ�#眗?ysF�Z�A;������p�3*�2�����1V��Ȇ�n��`����2����*��G��#�6���X��Qm
��9����9�c��K���l���p#&L[�N3�}��?j!*^X���8� S���H��q$���gۋ`uyl��tݾ��I�l�" ��UA<�g����'�Bz�,S+��G�����!�;@��??��#^c}������wi�n�����8-�=�V�s^�}_(�U͕"��gs9�iQ�ZSQ2xז�q�O�!3������a����rj��{��<�W��m�TEg��ɍ��t�]��+�ł�l:h�2Tf۶3�#�6.��L)��3�Y���9q��r���n��x�<X��!C&wLhuBϋ�H���g�5��N����Z<�����M�P6P�����	kt� bX�º�	��X��_��,!>�1��l):���mh�j�˟
鈦{��U���.@'u ��p��F冪�o]p��4��P�%p4�U(ʿ{�7D�ˠ��b��d�C�2�pĪ�m��oP|��q3O��Ң5ҵ�\(KG`���"�+�x*��qK�t�'�|�%��NK��T�@��!�I
AA�޹y�U�?��|$D�F�sK7>����F��|�509�k�(t3:�0걐GG i͞�)�F�u��SٮR)[��c1�g�5�s�+&s��r;{,Ƶ>�u6��~NG/ƞ�_M�f���`����E�| ��ތO�)7�2���P�068؀s���\����U��{G���a�eu�Hs�o�4�qg�9K�AU�mLw�9��F�o0�/����_37�{[`�[?�v�ʃ�g�G�궺t��k���I���n���M�p+-�3/yiS�#ש{X�S~~p�]89����=�;��A'k� ��fV�=�b�j
aV�>��1�c6���3����tٴ�Sm����2�2�2p���I�KLepl{�v��Cx�A��
VH�8]�J����+?)Je�������������f/KݠH4_�pA��\�(�fU&C�+��q�U �����:��$_�3͑�(}�I���ja�)1��r뷍v3� ���������g�ǿ��	�����hUƹ\��☮X��?����Z�����AJ��;�H�-yԉ�9�Em�T�O����w4;�����qi/zL��T,#�b8�V�+��c�ʩyVw�Yq�چE�����?�sXNQx6�+�����へ�mB�3�i���o ��g�/Ԍ��=t�8g�2�������j^Eu��Uw\*��pb��D<�i5z�i|��藮(D,��'0�;�l۸������,vשL�o;�Ҡ�v��-\c͉�O�8���9ҍ�j]��?8�N�17�O@�u(0�a
�	��2����À������y�d�A�.��)���1c��YӰ|L�Z�Al;���5���X����?�i�캮�ÿ*>�?�}tI�p�͎�Y�Z�[}��!p��σ�VW�C����!�چ�#^�Ap���*�0�ޭ��pT���Ԅ#�?B&6:��Z3�f^
|Р�4��8�1�Wk�b�Y��[�MgL��w�i1�8{�����V0��[ޮ+��|p�-W�\��X.'���)�c����S�JI���� A�c�ɠo*-�Ɠ^�c�6�l.ȥ�,���R�u��z�����S�����������F����~����g��o�Uc{���by��x�𺖟%�`1�#7!"`��A(P��xx"�Q��`%¡�J�k��[��͙a C��ƚ
�ݰj��Q�%>5�g��̒���s�L�Z��<Y(>��R�]���#"v��HzQ����$��Ke�E|�U�0\b�#���U>n�s�u���a&���UB	"��f"���w5e��N�z�q��X��%E5GZ"�
ĸ��rv���x썱�!B���v)�x�߶��.=/�!S�o�m�"��ݬRG�br��3��$�Q)[r��d�ͨ��zh;a�vNlT�~S����T)Q��w�j��K�(�^$��[�=��u/�5�o���f5�� ������7��^����{��g� ����߻���ġ�GK:�4�/M�l��6�n�12����W��vC�`�qȾ%"n>��I#U�茄{>��_�M���h�~`EEQ�dt�4a/{���c}�R��讋�r�7���ZgU
�7��8��hJ�)oT.,���X���Դ׿;$��������_b��o�ۗ��
�� 6
W	�����B�uPqS`��'��Q���v�_)d`񯇙2��o:��@!	��˥� ���v�
4H��H���cϫ�-�_zK����$�l�,`'��f��W�پ!>�ANO��b���>�v��PҜ3�w$'©X�w�zl�Ui��c���j���nX�b�,��1��Ϊ�t,{P��fL��h�pM
�Q�ޚ���범�YoKK{���Ҩ{J3�7�C��w(���?5�K�Ѧ��+���Tkk�X�?�R�J�l0շ��6�S��	^*7��_���.C|I��)B�)��,�:0q������+��Eݓ��þ1B#�#�K@Kf6�b,+bŁ��3��r8���S=�n��2tl]�r^
�r��1�0D#���V0�Ʈ�0}��O��eg3�I�������.M8KM����ULq��ǜ��^�8� �~8���(�0xd��1L�Ϋ䣟�s��+��L�)��bݎ�j�s"
Q�tV�tr�!�͐�*͸t\�VQ��5z�2�����8�m���;V?�Wn�= �=1�/��G͑��zq!�M���H˙f�%!��ѻ� �¤��[�R�6ѕ�t�)x�( <�'�~�}E#6�oeB$е�R-�t��QK�t�߇`ߦ[eƐ0��gEl0Z���%��� �Ê�'5'�S������B!��
d�3=��������Ȟ&�@̘1��(R.R��?�����>�z����Lпe���8