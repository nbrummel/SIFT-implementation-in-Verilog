module GaussianControl(

	);

endmodule