XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ǿ� #���_�������Y��VK!�51C}J,i�M����5L��^�j#�;"k+�2��5�/�-z�x(�.(�]K�
�RQQ#q���	O�{w����6�'e�rr��X�k�����S��El��wh��wjdb��h��M�ͧl�|Ĭ����<�jګg�ܢ�M��.���������5��ŋ��DH۫@�j@G�������A:F��,}���I�Vn-G>�n^U[�Hxi�ҟ��W�s��'h��z���G�����hz7��/ ���m&eM����c*��{)E�odjJi�*�]d���4O�m��P��m��ob�H*˙�� hXG����4�Rc��ky�\�"����R�A��$��*"�jzd��ۀ(�E��W��f��Qܕ�MV=Ju�ƽ�����E�`��F[�����f9�J� �9]�ơ8#�56b�òbȽ<���UDd0����}h?�V�OR��r��ע��KY&����*�	��!Rkh�.,a,Z蹳�:�����e�v8��v� -'�X2{�,S�Ӎ�5���|u?	����w�ҳ�6�md������q,�&'���:U��ު��k��y����Mo��0��<������R��[�J�tZ7��ps��ròq�rOYbD߀r�+�dWT�dZ�P|'cҡ��h��ި�ȾyN��5��Ů�z+*�Gy��=®6���N��k���:Oq��+���y-�
����V��,�%��yy�*�Yv �oxzD���i:XlxVHYEB    33cc     da0&���Z~��p��b��.�i)�)��[w�{���]y9׵���J޵r)�#���1�^�]HO���
�N��?��2L-q�� �@�TqZ����������<S"��f�o���g��'kN����3C�/��\�fw�wԇ^Q���?G-ꞡ���=	�c߁O�ݥ����uY���yGd�p�o�m��������-���8!`�|��[-���A����^"���B�Ц����&��}s�)����(\������rͤ����ovB�-��y�qVt�>��3�(4x��䐬y�4:��4yT�PI�Zˍ�WL��h⥐IlI�2���;d���NP�C��r�~~pӅ���,��g����
�葦�Y5i0FZ�pQ#8-tMk��\)��S��Z��4K�)��������ź��v�@}�MK�_���%�nr;T
е��D~]�qG֘bŚ�е�uhDVS�e�*b�a�!*�0ɯ���IA�w$`��4���{r#�,T�w�~eƥ&o8s����U��?Mx�DL,��$7.�~Њ�XC�H�(�����,�Bp�Q�$�J���ZѺ��Sڝ�K�W��:��+r��>�8\^z[z4'���>�[՘@#��mH0}�f)��C�at��޷���o�zQGM�r��$�����3+5Pq���Ȇh8Wp�,��i)�ϰa|��
�I����~n�y��&v%tK�U\`���Oq|Rw~�5�Y�Tܶɒ��ـ�b2��)~�����F&�u>�Χ�pl�C�<(W`��
�p�_gb����k�A���p�T̅�}����x��������ڌ�`�2���?x斔��{2?	�-�+����H.������M�a+�������?�������� ܄CG�y��_8����JQhD�&$� WU��Za(W�CtL���{�K���$ŵ��0+��坽F�I�d��p����vrF�g� }r;^�4M���$���C�{I���Jꎬ#�BIs����VF�*e�LK_R�hcu�ݖ�N-1��ٓ;��,Q��D�h$ͳ.�p�3�	i%U�	�ӊ	��H�C	,�>�!Zq��WA>ݦ�1�E���!U�͕�J���q,mJ%8�� �g�������Ge�]IwOABt��x���o���)�,��0�WB���v�cW� ��٥�$spמp�X�kB�޼1Y?g���p�%c�^��MG�i��yg/��� /��E"������A���r0A����a+�Er�i�9Y|~�'f	���P���d�/q4�
ɵ$4�O��`� ������I4&Nk�<�б�f_�ѿI�-=�o��2��n����[����9���v�=Xw�I����������5)!FKQT��}��0@��K��Zu �!O�bʠ�o�m,#W��0`酋�{a�(Ե���@ߵ��޶�hA 8|i8|>g{	bBi���۟9����%���ާ�u�L瓤��>�������4L�,�\��w�\fQ��|�1eK�2Y��ǲ�V�.״��J�Κ-�/��\���!���k^'�I�t�zrb���S=؍��91Ӛ�`�hAf�����E�qBK�����U\R�v��B��d'�~���b��%�r�sz���Ŏ���8�t@�J�/K�a���30u"��*�k�k�~F�C�'D�
}�!����8m*k��!Ж5�Ǭ�ᶡs��4/��_Æ@��a��j{q�"Z��t�ΏJ��,����$���O�,���h7���:�M��)��8~+M�b�<�����[$p�����&s9.������VgCR ��u��z=�*5e\�J�i�Rͣq}z�&�a���5�a��\���:�����0�=��Kw+H<�m�)ig����A�+���'�ۂ]�MUsV�z'_C�ͶKؾb�5�&-�08�5��������q�ࠝAF�_^0�������zPv{lڰc�E[s�|
�rocn7�����Ҥy���q"�b�ѣe����'O]f�\_���P $��`���3f�B�V6҃����}���[����.���]>�V�$�D�� ү�H�r��]�u��e�M�WW�afo���_U��ȵ�&��g`�$�$���������y�ӺeX��{��yum�e_m�W�o$��?CS��O]WM��75�+_b�B_"�7V��K��KH{����u�!���8Q�ε��M1k�����^Rb�$�}_\��&>a���'�?���Z��W5-)���/S��}��R����r���dN`s6�3��xq�)YZ�1��[��~We�5��-Σ� �� ���:�{G�!��C�jg_�qR��� 1�b�B�8�F�C0e�'����q�޽{�e~.�]0�!��ku(BU*߽�O�I��-���֩�A?ɫc�|�C��l��$�4�Yj�����&��L6r�8��y ��RD��C�[�/'�;u\����ߥTfI�C�Q�ܰ�8����@��3$N��4�_�hՉ	�U��td���h�a�b�I�]���h�����ʹ��sNzP)�� ��8��m/�i����J�����*���߀�,���BD�b�s!�^K2�SUoҹݳ4_E��0�5�8܇ׁ	Ֆa��K�t�hӾ�I�"����&K�7<�蘄��P{�foS}��'���RcDSt�g�_��\0��c �Q���
A_^�Fn��{���_x�@�N}0���V��!1h�pmv��u�b˽;oH�j�u��{�#$iN'�c���5V�Q=�5�U�����J��9� {u�Yl�j�]&�|9���ۦ����~G���\q�9>���sg-����?�w���)V����	��K�q}���{�P��t�5���qn��@�4d�J��d?�h��W���"
�B�p$���a7�K��Ja'ND��Ҝ-�nt(*J|.RO�1n�r?�K��g�\���6iy�.�\� �Ŧ�S_��P����(ل�e3��l������
�O��x��XZ��wQ��/Eg��}:��_K�-�U6V^-�`�r�%1ݕ�;5A�ub�L�vDF��
]��U�r�U��U���܄tXJ��"�6�
��Uy��>�(`[�ƆQ�����cWW5��Ɇ��zpT����E�"�_���E�Rd �"~b��W]}�?�	^����`��9��0t�8�xVj^�9�>0Q�MP�kD��"y�~[��ف��#��]ث
�~���� ����4���q;ݝ�,ӭ�L��	�_�:�޿ȹ!���3��)x�$��g��1��OrM���6D�Ya��ɂ�~���J��A��ʅҌ=��Y������E;P�� �tj��/�^ [�tk���C�^��1D;�5�IySt"�����%��E