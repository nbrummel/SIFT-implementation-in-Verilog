XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e׈��ɵw�N�[�C��PI�53�E���%di�P��[ 4W_G[T��\��)�K�U_���>ī��+Y�&ipo��?�A󈜆9dj��dց%�r/�س!{E5�Ք�d��í1�կ-N��;�K��Qr"�����b�B�V5�IT́��N�]O(A9��=���'Z�a�O`'U{���^�7�o6�	��R�v�ǀ	@>6|��T�?�ݡI��V=����sҚ�����f�>^�&p��v#��n)�k�Fc�����/f��+D~.���ӏ����,�AZ�-�U35�K4�ښk��:����竌/�\���G9I��+x�wb�y��Ѕ�L u y
��2�Ո���"p�IOV��|2�uE(��'��$�u�,��lI�.*n�
/�/y���O=�Y��/��3��־��<.�?�+��;>5%�����x^H��|�Q�r�.^���)�Q��L��}d`��:�D�9m�Xd�����Js	��h��������[��]ͷ�`c��2��f.���V�I�\,&�3��qv��E�s����w��d^dy&�t� I��`o%P��ن]~Q<
B��g���j�����d۬«���	m%gD;��M˿
m[�U�~宅{���~��5k��-�	%��~q�/���������}�tlAyf�?���z5i13[�R���#�
�q�����QD_�c5�p��UL{��U}[�J����$q��ai.D�� ��g�XlxVHYEB    3927     fc0v��]�,�޵�c2�������)�u�4����-[�.��>4"�U�F�<�.E)�Ts;�:z�a�"��E���<�Z1\���%I��MJQt>%ඎൗ����	�Wm�lȵ�S�8�)�=UV��4�H����泘g��Z���D�<8���0��Β��#�D�$X�|6�����nF���D
�����8�"�z�@��0�QY�ڠ����
�\o4�^4�g�xho
q#�z"'KJ[R�(SXUm0�鯨���B�k��Op����؉AQ v�|�ّ�CR������o�1}���w���yYqr�2�A���1�q������~��ᤊ|���j���Z�*�{�y�)�Z
K]�LdZ�5�e�R��W���6C�ֵSkbd�M��Ẁha�Em���0��
���f}�,���:i�@��_��y���-��}�M�����^����tp�1,��$�a8��>z���]߲��#P�s��,j�{/0}Q���n0
Z�&e�W��'�̻��~;.N�(�S��''~痲/ޤ�K����|��9*VaXs*?��LS���To��������S�|��	���L���)J������/��"����`dV��>'�;�?�B,|��ϸ��<W8`�)B�P\�Ҡ���Vu�u9(Eg�5i]�7����V��T����cO[f��NF�0�Zi@��2x��l6,i����X��|���D���������m��Q��V(�vmB3�Xr�F�ʎ������*dC�uh�x����>{y�L�U��g����U��a���\�"=��a�$}'�Wa���3����<�]I�g����{[�o�4�s��u[ȯ/Kef��tx�l%W��x7vm���T�Ӎ:	�����e���;���FD�V���"87�T��|���z�584��Gt�=2���=o��܎����+�mq���ق��`���u>�×=�Nw<Z�K�zi<q�s7�|/�U�4 ��E�uH앮M��ߞ��O��|���z.�n�3�4��:��)yu��9�Db4��[��\�1qok�k�3��ןP�O�ڰ@Ȭ�H����E>�����˥�m_��:�gHR1�*���P�B~^�/I�3K�y&����EE�x���|7�ʸ- �rNzx�a+^4�.��Z������	�����iT���4��Ƈ�<x�
�͔���Y��ͩ/y=�Q��5w��x6-[Џ�=9�^NE���μ�(���ֿ/��V*=Z�8"S�6��2��#}ȼ�60 ��aFѺX��`��}ʁ�
y�(���pMY?�rR�����F��塷�4���CMJ�0k��j����0/=3]�P������2�	nxe,pk/�!����(�Rc3@��<Df��L�������3o7]~����xi��:u@�C�?�&, ES��3���^�U�|�:��W�T T�v"]�rE���3���3q�mPr�0�o����B�fW��j<�^�6��Q78
�����9
�FP�-�V]��^�%���`'=
M�IQ�W3�X�gkFn[�X��NphO�a:� =��wy_�.�jQ1`���溅������6�����ܖ���MK�e�ZY��L�]�2ц�΅�P;��*0ҩ�O9��G+���Y����7$��z<��n����/���3��a�ri0��E:�% �UW���J��͆�;s��k�����H�3�y.xB����h�v>'W�"~��}�Q��|�XsX��mL��'BK$�F��6=z��X}�~�{�B퍹��F�XY�=ZC��*�t�g��6e����8�>oF	��Ƞ6 9XNEq�52�p`�a'$��M3�]�{ԩb�ϰ�����(��_����� ц�(q�I�D�N G�����KS��	di�S!�*G�ZY��WY�1+�%������U�9��O(��=�A�����)|ݙ}䳄z.S��Z����=��J�)A�<��Ǒ��&)�o���j�{=�Ľ��y�[v�Gmz���e(oT/�@o�k�,Ŕհ5O��M�����F|�h��-����l�,q�s���:T�Y*�������HQ�" Q(g��$�["�/O!/Vø���j�,��}���M	���|ᢿus�Y>B�0�+�q��U<�u�3ӑ'�`��*
�x�U*B��k����_xd��}=<�ں9�'�	�ꏗ5F��j%&���'�����%*���r�>����:�9�e�O�םO�F�r��-ag��R�2a�H>{�i�=�zG�0�~��~	�����1�e�[D-S��F����_ �1��骈 {�9I�����X�Db>!�V&��S]L�7���b��Xs��(��ov���i �Aa-��9m��N�L�)��}��-�)x�N�T���b0.����?)1���>[Þ���zܳ!�i� s��K�A�zkx����]x���ܕ�א'�/�
Lh��U�J���ѭ�lU@�8麧zT��%�6�U�e�溌�� �`zq5_]�;T)�Ku?���d�0NOt���d�ƚ
�:��9��X��qa-I�EZ�b�i��ħ#�C)�v+vٚ���zm1}f����L�MT�9MbS���{V�q*H�"�X���u�o-�++~��#���Һ'�e�Q�dB���\�<����k֐B��;`�Ojd��d¤�T{��/܍s]��x�7>mr8"�	�yU���pyNb��F�x���I=O�m����oG��iP�<���k��d�&}Xg�F��I/-S)�S���X��/ȉ��&O�_����4���[Q� ���p���,7nh���Zڞ���R��+1`����뻬bQw�QiM��vB���i���و�+��C!��uwK\[�ޢ�y��@�� �����sW���[������������l`��R:2\�(��u�� G{�[����-�j�jV�v]+�0�6T�Z��b�@�9G���J,�"u���T��j�k�'�iV����˔��d�ۿ7��mr|�_a�ݦ���ڡ#0�'�4b���XTM:7D�:������̮5H�Oh����� F�7C�B�
ラ�D9E��y�m�{�%���7�� ��|ͶvA����X����,�u9�c3]n��Y�D�� ��~�:ID~�wQA4ڭ���Q���j|ê�W�b��Ͱ
���/�A��g'%�j����¹ڼj��m.����;� ��XT��T�:
L��?�rE�����nT%r�J~YntN�8竕�ꠢ���v�:V��aq�q���ލk�so%��}��4Cf}�rs3}��m-�L��漦�t1��`��>H+(~#=9��Y��!�2�`X��crx�T/�"�H$�ꆤ>"s�dL��Y�5/�n�ԏ��V)V�~�C�4#����]��k��?����s5��g�"+����Y��	ք��|���x�M�d�n���#�F�F���cU߆QQ�f��@��A�n�?
�G-̅
�f5Hγ�N���-��[�Z�9���[����U�!�A�"��@�>Q�Sh'�p�7Xܧ9:b�
�#0�畢K��A�T/���UL�o˽Mby�a�Lчw��÷1�SX^1�Z3�/3���Q�s�n 5Y�J6]�訁%�,�&�6Be����%��������[�ek�9!Q�`X$�`��٭i��&R(f��-fm�v	b�(bW@F�5U��`�K*8���^\PF��}]�>��'�F7��g�_??~CV�o�eU��\�Nl���w�d��D%U�*���ٷo��u�i���a	+^�.�֜n�8�6jR4ʑ��޷=��n�=��oA`��MV�ҕ�,�YS\'���l���`�A�H�ޟ�;
3�Ss�k`R0��
� ��uS��T�Е��+�J�/���"�w.<9\�Y�&2>J���h���]O�JH�(�M���N���!�ߟeW92ؚ