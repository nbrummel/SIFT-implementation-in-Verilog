XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G�vHUZ�]u�|`#8�aŭL��NB�>��V��]�&E�+x�0�2����ק�+3�q�*/���ȷ���f�_AS=_�8`��C�4��&6�� :���H�t��S��>-	%�q�����n��CA�dc���?J��j����w`��������!�ղS�-3��[}�2�N� �*i��9��TB�If�.,τ0��s�Ύ�0 �1��Ƚ��ub�/}�N0W��ԯ�U�Ś|@ԠV�!��2��a�nʓ��shޢ�J�RD}�K~/�d�X�g����Q��w��ۛ��z�7�E��A���><]�TϜap���"B|F��;)��\���3ݔ�Jo-B�2KIde��F�x����P�H����7��B̓�O��v��ui�$t�k�P��Êu\.w�(��_{���s|�clJ���[h:3�>��H{����P��Sq=��Y���&i��~7tr���c^$��йX�	�f�W��#��P�CR���(N�gZc����˦]=����"ƣm�g�iׯ��qc�Y��qhY�SƮ=�|׬H;� 
�1�}h�~ͻC��#��rtf+d�Z<c�L[���xp�sr-uX��x�T�X�3���<z3AS,��4��8�U��&I@nk2<�+��q�-�29�I��2�O;�;j���TX���'��SDj��^"� ]�6��c
Ӎ��=^kX��Bcb��8M�H��]7�})�q�*%�EE&�c#"�ɻ�&}�Zx��b�Ԏy*�XlxVHYEB    1802     830%N��-.�J�%�R�w�}a������4�\����W<7��B�@�ēmA�4�a�iJA��D��#u�ID��2��\������D��'DK]eؾLR��f^t+?$��Q��Ei���"Y�yJºk�r�y(f�BЮ�7�lʋ���r�k{��\/�l���$ľ��^~*]D�l*��h;����f�����W�f��PK�Ek����Z~�,�m��Cl$��Y?.�{/�':��;��qG�����Q	��k�R���̻U5 ܫ�c2~D�@羞�|b�}�J c6�h:�@u����7.���F���<ѐ{���;t_\����̺���\�3�M� 1����;S$���Z���qT�V�8@.I��V0��`���[�ڻN=%�^���:/Ĺh)��@!ac�6��E��V-bq�$
����}��#W����
�k����	}ה�{�g���g	f����Q3w���C�D�E��2a���0Gt���k�Q�nv�Q�>�)}CcP�Kw{T�!�t6���tȕ��~<�X�2��V���=)h�!��Y
�$��N^64�ż��o�ɗ���2�TN�R�l�q;����U�؅�uI��U7$�:q���˿)��h���ߝ�$DS������,��a�g8cL�.�7P����6&7bs"�i-�l��J>4ρ>��BE�׉H�?Ғ��V�s��Ei���a%?��G,'�HV��*�D}H?��"k�*�\e�H�Q�;>���ˁ5�h4���Z�#D,*�&ߩ7����3�B�s���Fh�@����mb6Hs��Gfrpu�㾑�R�	��f_���e{k�㙿'=���<P����% ����Ғ s,��m�Tm&�`��F��Mv�N�0�&�[.�qki-N[q�+���m@ԫ�R$��j�.C0#�:�ձ�����e5
oimF���^��T�����S"��ɃL4��=���x��F}M`��U�3�|hJ�� �Vh�i4�hz�j�����]�_N���fS�N�bd��O�|Z�vΐ�y�x��t ���j�<�6Q:U�l���tk��E��v��x�8���Yg⧞bIVO���(p��a��4��t&�D=Øu��F�~������jJ͛*��|����%h� b����}�H4aBpNg�C��&�~6��Q�_��oZ���\�b������V�3���0��f��Ϩ+#�����G�$앬���d�������NE�^5;ȑD���`��~�e�A����B�MbF4�調�7���Ugl�nPB>s�m�-��VX�Ş*�"�C���,���%4�)O�P�y�4c�a�J)J�������U�}�0����L�;\����*����F�Z.xbf*|�^�7�k&��D�O�l
�hm�Ls>�"�� 3?SsA�/㾨?S�{̸UL�M���+��QƸS-9J�ѵ�%6�\�:l��Sw�'�	��s�����f ��@������¾ �L9�1?��~�������� 5���R�q�R���?P_F1�S�� ]	����V�+��d�F8����3�ԌwA]��k<�d��(�_���t�䒡R�Ƕam��c���i�S�mBD}�D�Y��7v#��L����5!��1���}���1�h�x��eKᥰ�pbc)e�� ����y��cvI���f��o�d�"��H�e""k�PC�����Y�NYuw�����n��[�P����ԵR���wu�����Y�`�/#/�����.R'�+}�^��ě�� �ה�^��`�c�8�P��;,Sƻ����ɒ}uZm+B�D�w�W%�<8O����9�p[X%%��~,/ �Th�f�~8ݧ
��מ,���0��v�A����r�]�T��9r[�)�^4z����GX�p��Ԯ�����{�����cx΀��X	�;��sЋj�P�)E
�G����	Q$|�^��PgG�:�N���:kxD�-5A����RG�� g�U�Lu	!<��ʰ�BT��%�9�h'�|[N ��MJ�"�Gt{�ev�i�IZ��ܹQ�
�@�P���F�v� �M��q