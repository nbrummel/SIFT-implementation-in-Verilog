XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���/�F���cT]D��p���P)RE���N�}f��:*wLf�H9�ͳ@�
p��d(DZPjxr!��=�jW�2�2����G����D���Pjp���.�R�����=�Z�!�H?A���!��*'�eh,��T`�����>��lRӏ���b���"��d��MfnEq�����4��d�VH1�����o�:u=�j�3�k�eq�����Y��>�> �8��ɢ��UTأ��m���]������AMC������3�¾��R�ЩL��h�WI*���+�^��舩�fr�\�n.p�ؑ�7	߂ǹ}�׊c|Wf�K���V��`��v�qiL&�ru��;GɽM-�B���o���紾�(<�XѽU�n�.*)��L��)�Y�QS�۫�vA�zK~��>^X\��'.�\ǆ"�B-�����N}/m]�����l����m.�p|:�?�]�����C7�v	uT�H쮕8�L�<�А8#��v��|e�K��n<M�v� �;�y+�[8���/Q� ��t��Q2#���!����&e�'�>�0ݢG����BI·A�S�V��y7�� �������p�72D�4� ��U�z�ab�U�;	G��F���"B%0h �N��p��3�&{�=�~Ȭ���羍G.Y��غ�\��D{�3/�_^L�K�K;������5F�K�r��Ϟ��kN�*�DB�[�����:��0��%��Y��]�@p2��y	��p�XlxVHYEB    17c1     810���#3��=u��̋]�h,���Y�
R N�u��m$tMSȢ�I甶;,�./K;!��o��2�+X�8�����0�Qxc#	�-��6���ˎ797�#� 3	�"�a'���d5� �HU{��2�����1�ؑ>��GH���EJ.�E���]c��E�=�mծ�����Qw�0l�2`P\�̬ek���M7��j4Oo�<u��1���_j�������bkM���R���Oh�U×� OT_ ��\�3��2p0�ѧ���j�D�K]���L�TR�|�=��┾	v'��<BAV�~���;qB}�M��90������| �����c=<�����bL}ț}a���E�ni�$=�O:L�gp�F���F��+�Q�+�a����E8C\�<������i���<,i���J�ً��5Sا$-��_}|��ŵe%�V��%ȕ��W�ܫe��y�F4I�al�Q~��wk�A���2	�S�zl�Qv*�ƫg���>�y:
��KgԱ?�����j�Y]i_;N�D���y�>������2cW�Zz��6*O�7j��<��a�� ���^)�ڣI�➉4�����cT�̵�yi��Ipc�I�[J�W��ܩ���x�=�6�5_��
]�=tʱ��q��{2���|G�͛M?�D��O��k�
�i�cs���/��E�0��[R���>n��
 �������O���e�;!Vf��ug	�ǎIT��! �����Y��Ni������u����׷	��p�>�p��7e�I~��iř��_GȚ	).���%�u�q�;�����������=�YA�/Ƌ�aUzB��ⵜ0A'�i�?�`���	AѴ��W�Gv=��=�\�r\��F�7�`���~�����
B��SG�	�F"�N�p���챽�lP�u�ދZ��P ���`=�ʋ��I�{��oq��~9(��o�ڮ���oZ���J��a��7y�uf���sC���Y����vU�CY�f�����C�ӡ
L0�+�M/W�r����]x٫�%pE؍���i.d����8k`��P���3�+{l�Ҍ8�'�򙹋�[�He���5��bӳ(��|�tSjn�/~]g�$��}�ǹ͛��)����ƪ�a�1eܫ�c���D6�,�B��p6'V�1c߈_��]�P��#���D���Cz��p�a0J����Ek�g��NɄ�����ڣ�|�N�W���IK� �U�I~1���n�V�'b�j��b�Z�?�I���M	���
�h�K���1R�jPL~{x�v�_Ȳ(�qj����Y��=�Ņ�B��&uCQ����i��s�d--T���K�V$��2	��&�e�e1^�_4O�1'$_�V�����&_5�2}����5�}��[�ex)����턳����T�O�p�"�_�P�}���W��i%�o�3+�l���L�YU<$"�{K�y)��q�3��HA���<ub�Ex��J����n��T'CR��Q$��tm��v�w�����E5���[��;׉D�QDDS��@��*zH;���t�߁T�_��v��HfI
��ݬ�O�Tnp�������T�����A�tL�f��:Fد�āטw�������=�%GHplHde�kr��⹢Sؙ�﹢��`ߢ��V Ȋ�B����ሼ����F�	;��(���g�i���Ir�l�j�s�l��]��ϣM�qx*c���;p�'�����?��3/E�~++3�������*���$���i�[��g��:�.���s#��Me�4��?ا���4�&KU��o^���{.�1���X�~��&.�|����4�}����ۍ�Z[���m��>�}�N�����Yͼ�Q���~�n8��P�w�Y"O|.q#�H�	j�U����dt`u�[�ҹ�&+�0�Z)�U�bS�B�i�Сذ�@戲U)��c0��T��#��p1�B�	���e&���RYI�*��(��� 
+��H-j����_��
�e3�, Vk���1��X%8�Re�7`