XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(�Om�~m��Hcq��$c�%���I���5��as���?�^3a^��"�ĺР���Eʭ|�m!���?��.E����"���4P$LH'�f}B����K�
,iK�i��ߐ`����]�=���B���L�ٱ�#�'��Ӱ,������P���F�8���?vnT�����G+�w��˱�b�塀sV��3���g[�5����7 ��U��{u��>��� �s�| ���?�3����,�w�0!�a �)�۲7�Y����V?�+}�o��G8[�A-3z5�Z	��YK�ܕY�i0� �
�V�&x�T�R��e����s-���XcC�*`� $7^��+��q�~!�z-�^�q�e]�}���u�@�t�k�2D���=�>��@�wPl�*��k�v������DI��ug����t{x'{FK���E͛o�y�/ �./�|~B �<$Q'�㸟��[��!]��ë�Fh��AD��믎[~�)@����.ΰ*��޲�����x�h�ŵ�$�p��C0���RL#K�����O����s�h�����Y⍪���m�!^�kExCO�8��}i-F@�|�59_�"8Ō
#�		��̤�����"����@��x���	~TqI��Ҍ�R��-u����2M,�76J=�Ma|�����w����oǷ� C��N.�B��L0b���L�q�j�(��ߋiP�h����"!���3�ȵ�q<_���w�cQ��*aXlxVHYEB    66ed    1670��S ����1�����x��mP�z3���{�c��K��y�>8���<�F
������JQ�~� ��q���W�J#
����R����b?�[x�ެ����Cb�X� �ܥ?QK[M�v`�<�x+Z�)hn���B��zP姚;h��/K8��l�	h�p�xK�t�W}u�� V2���Z�>�J�zZR���}K���m���տ��Te�#2��u�征���_�淖X�T?QiM�b�3��8�Ս�����`u�����I��mZ�5�4x�O���BKRƵ��T��g3�5�{����.O#��iE3Sq?�v��d��^�U�>�~�w{D_P�d��:�LG�&�Ci�@�a���������[w���H�	�@�������oӼ�N6����#�V���̏����z��wХ£w����n�C�R2K����<@�^����c�Q���j�`�A������Ks� ��o ����/Ɣ�#�+u�zn	d���W��cj��3�qFf���⟩��Y";�S���{�ϧ�nRP*�$$x���z��7��q�u�nw�v�,�X��܇�a�Pߒ��P�85��sCƢ����
)�m���'�Ӱ�ߓ��w	��e�Y��2��60��IX��`�������fv���o�h
)i�1l-���N���OX�e��R;�3��Zef��:'�q�Q�
�tJU[��P,�&|���'aJ;���	�εH��6�1� ,�7q��M<���2F���������km#�`cKk�2���b�RW-ɘ��;'q����!�h�l:�}`�*�J�[l&)��� ����/��xw�1�<i¨�?h��e����<�?oH[�Wx����|���7���}\pvY[��9�G�d�1��!'�d�
����^��;B�h����,�]mE�T�uz��A�[:�+�
8�Ɉ_U��@I;�(���5��A��^�>�
�;XN'f�5��a���Ե�X��#6@�h\8���U�6I8L#be�Kȼ�����X'	;�7v*��]S�>zLZ-�!c� []$W��|��O�g�\�x�҆��{�=���l���)�Ȋ���Y�S#�[�y=�����*���8�k�~��X�$��(�&/���<��g	Y�2z0BhT������v��6w��ȓ>8/��2~��-B?옩���q��q���m�u��_��"�1���J�F9�,���t�r�]�7���@=�qpp���t*eEA;�$����"q�!Q�(�@:�x������\�
Ü�A}�љ��[�{Ŭ�ڼMA�׉�9�ezGҏ��_����
��O�Re(2~�	)��+T��Zg�\ ��n�[�#��^����g��L:̋��LTKƆz>+?�5�3���QJ�b����A�a'̖[��P������hU1�9�H��Wޞ��]�@_@�qVF�K��O��T��*��&�Ah�����$me7:-�$1D�S֨�2����v��7fV<RE��?�hOj��=Z���ƽi�K��4w�RA0#�ٛ��^�����}��8CG��j�����+%CȷX0��R[�Q8�01�����;�W�յ%��c6��"z�҄�H���̲�(L��4-����	�����Z�7%�>ko�!Hú����S&*D;z�<˔�tr��/Fl��xu�J����q��-4�j�L��b�ϗڏS�^n&*L���{���Ud/�ՑB��1��DH�.^�y:t������;\�q�ja��(p�3`D%�LS�w��@���D|25�WN����~z������� ��˷Q5�u��n�)/���޺�s�'�x@e��M�s�\�O�_��AS��)av��8 ^����Fc�rB�]G}o�������K�?�>�Z4��R�	�Ȕ�.� \����F ���>����o��s�K>�3H����,�c)f��v��������1�X;��%��F����3}e���_��y�d9��D��P�%��>�U�ͧ?�[�d];�azו�ڊ[�Ĉ�S���!��/�uJs�i�eJ�9�Tw]-���?���
?;���`Hm`��n�z���,$ ���L�ZQg��$�@�qKԊ�d`/���l��tY22�l1ƞ���0��h�?��SĉP]��V��O$��f�M�k��P3)�p�����X��k�x�IaO`�Tz�z`�邨�Scn�$]-�@9w����22�@�ge��,�.f$��� ��ZJ��Nh�bIOE{~��Α;�r�_@���=U';*���js+c�A� rn��x#�����N�n���F��
Qi|'����~�s �sӭ���+�5�j�B窌�)�L�Ŏ.:4�x� �9;@f����:�G��g�QsAVn+a�"@բ���ElǓ?��'8��G��­9G-�%�0�%�&�����^���Vl�Ԩ���{��F�8W�Eҧ�Wj�C_��l�@��4/HU�ǧ������f� ��zR��[��ҭDT��^^�@�O+}�����Ay�G���w�oW�]��c���2_�sP�L�{�4�̦t`	[Oe�:I��iv[�� ��bЊ��36�r���$FkR�����* � ��@p�`!������Q�Q�a�P�qc"
���48O�����?6E���e׵ b�.����"J�qw��:.�В���j8�T�T�T}q��8r��0��r@}�D(e]]:C�� �-5�n��Q��oV*���sv��j5J#�w�t���Y����DX�t:��2
x[�+y�9��yK'�����y0��l��2/I"�[��r�Uxe���8S��$!vX%�{^}x��*Æn�S�+�"|;!�u�bZ�ry?B���Q\]���*F�f�J�u���,֯|GW�� NN���e���������W1�d*Y����~c���@��P���/��e��s��	�,
`樄n�O~jR���Ys,8�iM#��9��q�$@��FK�)�/��8�f��{��7T���*����`�a�����S������s��zKR�(����s�J̜mՀ�cH�M��c����ɶx����4�
�&FM8��,�2�Aϕ�_(k^�.cح��;��<��
;ă�{�J��8�<�J=�*�X�SmG��y}꣝��\�Qo�%sF�@�cj���S%��\���̘>��(`�M�k�i�rC�.���]A?`�$2¶�d���ڣx�y*܌�AYԓ��م6W� r������o>6ڿ��L�����y����G��ٮ_��-,?,P�4��7z��Z�R��ܕ�`�-�@���QE�v�t�'�a5���?J`��������+�*��`&�w��S��mia�ңcZ>y���/r/�#�'��?��2�Ds�����27�nIۣ)����s;5T��WPL�T������P��E��&�Yp�d�	,h�t�e�@�-ZƏ1P7����,�v_F;纐eđ�K{5����6�πЖ��6�h��)|�'���i�+M��ʬ�LX�*���?����������(�UE}�R�k�`�S���:�A�+?ޝH���úةU�R�	�-��T(�R�"Jv�jR*ى�ö��5cE�?|>���t�Qs����OD�q���t4�@ g���=5�O�HsE�Kn�>�*��Jɒ̩��l�(�"�v
q`���ń|���������Ia�)4�|�p�;�Q����US�40yH�ؾ�)n�ن�Vm��A��P��V����"��s�A�D0n,a�RiM|���il�ž�L��
�x�����'���iQ��dD�\�R�N���%w7v�D� �-F��h,\�U���&pDy����+�c�E���@��;̳w�j��g�fv+�얿��B��A����R��K����\���p��S�'�q�_ib���x�
k*�[��q��m�.���6��V6e�\�mO3�B�b��/��%ĉΙZ�O� 7<A��c�!JL�J���N�S�ޣ�U~6�3L��|�����X�/O }��4/�&>�� ��0��
�c�������h��˯�M��8��SD�
+{�6i�u�V���D_4́��1�FAC���h�@�H���a�
t(-Z9���p�Ip��k0a�)3M�۳EH��Gb���DHL4����;cK[�7�	�/鈩����		՝�=�b�q��W�b���Yӱ�ir{��=ձ�ڹ�uyΟ��m�k�⚬�g�h �ZW�B�����o�.K�s!=�7Qa0��V��e#rx��^L�J��e�f*:��k����؇ׅؔqG����ѭ���>|�v��M�|�Q�)e���P�q����|pf�}i�iw�G��<����zo,į!���_����_����G��1�+�,�Ȩ�� m�Us;O�ʽ!v��3���h�[r��,�\
8)���4�a2Yj�����/��w`t@����{���>�Ql�4�|�p�L��1�%�ҵj�ky3���l6��������E� �-u��~A�I���C���/F�7��l	^8�^@��Dͱ�|"s:�W���1�ra���c����u��Nk���	�%pY&�.w�d嬬�����z���.��E�(t�hg]�pԣ3�).��2��4�|"�C�]/dm���\�<<9�4E3��.xQ}V�3^β���LRA�j�Y�O�fl孻Ɍ��M�B�m��L���%��	Y�&5|Eo�=�Vk��װ4�(��S���;�!�qZ>�u�Y��$7�ݤ���u�݂�x Bu��_���/~׏�K��o8����U�B��	�&zk;\�g��
��6]��W�9�ȴ�Dz,_���aXGſ��#�ˍ��Ľ�֫(��M�DuZ��b$�7w�\f�$)q}+ӖH�7�T��V䚋h�;<�d ���G�r�u7t���C<QM�h���5 ���6��5��k��D��2�׿����R=��g�ǅ��!z(
߃�95l�N�K��rp���qi���&�Z���J�ŭ$3�ߕ����i��I���6&$����m�PI�m�{	��䈈
�!�D>͙L��88rڎ,fʡHL�@sиJ%�[5㢸50�vN�O��"��LĭQ�����ݤφ����| ��0�)�>�#�鑻�!\���U���0�jV�S��؍c͹Ӿ����f�n�D��jt����v��!�f�؉M����	�`0q�W2�9�1xs}j��@~/m�k�@�����9DX���N0�8���~b�W�vu~�h�g9�����@�7��-�g��h���"�9t���IV��0��S��ڝslW�ۑ�`b�����AC��1��=w�w[RQ�<��o�
3/e�x�q^�Y�ЅJ-~�sCW��o;�5a�},�ǃ�R_�YP%�Iu����ὌL�3c�t��=xp���x�|݈�v.|����������;Y}N���U!�ף�6�.��Tg=��P��s���������8��T-]�pB-7v�5��~�[5����q�]�L�l=�S(����ʸ����Rqe��y$��G�(�)���*���j����}����]y�6#��QG~?����'k��7����ge�����