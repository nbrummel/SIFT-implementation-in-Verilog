XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���8�'$�USyLQ�Z?�����0rC�J����J��Wj�=�2����]�W}Fbh��,WR����������J��uD���$��T��!��uL��Y7ב}	�<+6�S�z��M��~��w�AE����i�F�<�F���)��%�	����ʍ#S0>w�ξj���b�ߑ�-}l*\ޅ)m3:�%l��<�Ĕ�P�M��
���Nc7���[V!/o�����&�u��T�7�n?�h�KTA�hl�rw�Z���D��c��eD��)��E�Ln�\Y�/b�(Yf��?��^
�_�G������v�Ʀ��;��~:؆u��jU0Q�r's ��/&�#vSS�I�G5���&J����5^ȓ=ʊ΂���,]���d��h����2�.��-+๗���tj���[_�X��D���u<<����E��r�� H�&W��\k,��D��m#�j)+R7���\5��(p@��_��{�ҭ�	����r�����H�c	�އ�O�=.�Y�:�$#S4�jFİ3n�H.�&�*Lh4QU�������7�ԚP"���^<��{O>�3�o���;�5��#fM����nmC�iL���/�"���(rՒ�����<�Y���z
C���'C��DX�,���iH;VK�T����3���������Æ����[����0��`N��s��{�f��������d�F��c�A�c S�d�I��V.��m Hт�!��XlxVHYEB    9efe    1be0�4����ͫ��������E�@oV�����IuXD.T� ��.��y�+���_��uB����9���e��<�V	�V$�o�!�őNK|��ԃ]��7�ŅT��H�(}M���ҢTt~]�1o�&��4C[�b:6�����:��&�C]�:��R�0���=��+�n'BVDNb[Ř7cR�;���1|���|���	W����o�n�U��w8�������HG��m%�$ka��A�eH���q�J�����m�&�PN��#د���{r&�b�>�h����5�O8,��'`���"����5N8N ��7埓����~fa!��q%JL��� �Q��&ǐ']����eF�ܙI����z�T1��
;![�O)q,���{�IE�R���o�hU�8������KBI3��+�K\!Ӗ�TU�zB7M ǩ�T&ʕ?n�)|�Y|��]?aO�?�
���O��٢�*��ŁΏ��j9_�C/u���O�������6q��p�53��b`�e� }J;�V�*ek�P�E�����̓F8Pl�#����s�̉��N��h��[`�>�:��u��"���ݝۡ2_ h@B�+���Ҩ�AG���ne��,bh�qi��I-�ҝ�^�?���!�$i���J�l}�86��^ӯ�%�c�m7�s�>΂�Y����9D��`qO񌻎���s��X�C��ɺT�'�(�r΀%�WC�-���Mg��ڊ!\���J"O	�
XH��4�
^Ŧ�� �<��,�(��`9�j�'�Y
��>�*��h��7�ղJ8��Șv�\���/�g�Ȋv>��^_��PѨT\�p�{E��}�ΪNT�$s��=|!fny�݉���z��Ѓ��Z��+��s��|�tai/��|�X6DE�.�	��~8�����cJ\�RF�/	�$���A�:;Lm�n m;JE�%ޤk��|��D�ˎ6��Q��{dtn�cr��c�$mݬ��l�Mq8@����:ju����S{Dp�o;<�!�� JLd ��8�tLb�t��O�(�'�o~��N%0@��b'��f�|K��G<����ӎ���p��Wh�������Qh�C���r�]�G:C��l���
��Uƙ��x��oN�լrb.lN� +���*�Gg�_&�~���8f����D����g%*��G��<G��J,U���W۹�$���ʷ
���Py���1�ѱ!��.J�{�6b+��o[N��ʅ��C��PR_�;��f�D�(2�0��{�,��f�6#	��%�6CR �=��ЭeM���N�����Z��
�(��SdqVoݐ�����\�$v9mc�lv%�U��5��j��M��tPD�@���ȜXϼ�!�j�zIHй��󀺓]��Z��Ad���LK��y����f�UI�S@0��ָ�^�X�6e/a��+Cլ4���C�g[1ڟ��*���<���rta���<��*��5U_��Y�^!���f�/P=<5�%�Ig���x��`ۛ��he/+a�͎�2�q���յ�Qd:U�.^�xW?����y�G@筥;�OR������0A�-y/,'9� ��AŰ�\�� v���|V����91S��r]Nր�֣>Z�j�+�v�$�I&��O������JC�q���#�D2�� ��d���>f:KԚߥ�Y$��5�x��s�ŦR����6Z�^����q�ʢ�H���n��:���~�Xw�!��q�T�{9��|�V�k��z��k� ��A�g�r�l�־��`��0X�`�(�&Ή�3U�5��r��(��C�������gxEK�
�hMW%-��`�#����<��u����l�&�bt�1� ��J�]\f��T�TH�C�9�F/� }pK(�����G�^2���c	{���W�	6�DT�!�j��
��	���Tq���H� I|��UO`�7� �X�t��
���l��D��>�H-��ʹ΍��H���>�~Մ��(�؄���� �a@�1sI~�Cn+A7r�	��k��]ʾ��2350'����QR�*6��MrOF�J�)�;u���OQ�����f�މ��(���h�9�W�L?�\�y*o����1�zS���YA/bH���o~��Z. 2�	��V�Ѽ���0S˄a 0�����P�h�x����@�N-wC���wڤ�7K7�l?/�h<K�,ɁBu%���7�3z��݈C�"N��LZ�����:��Qܑ�C�����r_��ܝ�_1*԰�����d�D5��:׬����	+!\�����=yL�����룀��C1����1���cp{"����z#�E�j6��D1i��?�P�t7�_��|�|����?<3\�T_���~�E,�UN��� �5�=�u��T��Rz�ƽ�|�4eF�tM���{��E	y��N߮,���O
��\�h�j1�b�-��j
*��-��@B�z��Az���� .7O/A8Yj��}m�v\@�N9�):�x7�q�n͡��X�eC4��ڦ�� ��eQ�%E��l)3�Q��y'�u�4��x������n���ݙTπ��"N{U-��횔9:ၭ��K���.�d�&)V��Ҟ�$�h�xoo�5&Sy�w�Pע�5Ea�ۋ5
�$���1u�L��;�|�ÎȵcΪO�1�M޷�}8<B'���Π�][u�?g���m]��U}�/��(V^�1����ɽ��N��WV�$*P!�h����rPWoo�T9�XJ�x��zм�&�?,
�85/�P�r@����>�hg[!��gC���V�pR��šݴ9;wx���p��%P�b�>,�(��l�+��j#������ph\��0��;1��w�T�+�֌|C:��M!,D7��p��0�l�\��1�^�.i�EH�!����LG�jD#lT��G��r�ߤ7Q�F��|FCI?@
�,<o·�-��5���@��n���k����E�G+ =�b���Ơ=#{��b��p�]�0B��?.��\%�)�R1$�
�)��;(��f����{� ~��[6�Mͷ�S/�΄{WE��8��,m��ÚA�='�&�|o:�p�&����``���et�ѳ�9d�m;���R�X:�@�(���y��F�?x�li������-z쨾��L勵����XZ�O��v���ҁ��n�z%��o�P��΃�������jGF�64��TƲ�⋢A�G��=Ɣ#��kn��9�������f��+�$O�Lc��@�T*�2.-��$1vF�F�R�[�����ާ�	QS,P�щ�%�c8b���+�;�`yդ�-ɖr=DIb�<�o� �)�A��I�(є�vL����Ɛ�O��J&���{��@K�q��#�)T7�0AX@�Oz�[�_xk��u�T���#�O��)�/��i�-B=y��vP��I>T��>���&�{��|���)�z������9��p3x�%ݱ���D��et �l���%�����^/p�08IѴ��W	��nf�_�HF�JBU�f���qu76iS)��{,T������O�l�ز
-�VEAwv���>������H�E2@
	A��@a1r"=�d�H��<�����T��q�6���Q�����\4�Ϳ�ѝ�n����#e��g�s;�$+j{�N�Rk{>R��t��?��mJՌ�8ݞ�-c6����g
�*).������=����W/�C&+9I���$���MBC�Ȁ����_��o�9��������������ZE�l'�kQZ�����f�����s�Ĳ)�q��1E�bi$�}k������*yjQ8�� N>��`jUI�"!|X�Č�����l��-xQ Ǩ'�wZ�I�ʂ�#�>�%wDxg�̀=�{2��(��>���Ǚ!�N΅�Ƃ&9�]��NX�$�ƿ���ϝ'hvW]�ǛX���SPDc�����*?u�r�e���[���5Ϥ�h[�Q;�@��|�drZ��Q��x����٥��0�>��L��);#�{�l�̙��o�?� �X���V�C9�9�VёkB�D�w�օ���4�=��Qh�I�R<eM�j���vT���<F
I��1JW�޸?ͪ��E��[P<��,x���$T�R!0��O����u�r���uچn��c�PW�����#���ݒ�yJ��3�k���:d�ZK'&�E��_��ӌb����⡋�J����3v5��&>l�M
��w�je�#s>,͑:ȁ$���p�y\Rvq����C,�S�10l�س��߀PL̡Nq�߆`şN+!�;;����.����M'�g� ��}(�4g�2@�C�䏲C[/6��S�"|A����G��-��,�>�)	�kW����sE����bfyp���65d�ٰ�%���S�A:�.=��NPv�\��˓�˄��"$dF�9a���Ƌ�9��h�9��m�$���Vk�}�wE\;�M'Y�Ov5�;%'�[B��afH���P���GE*M���7jQ�.I�j�C�H�̄QCC������"��`���B��F��n����<U���eB�C��f����N�f���_hO}���<|:���n]�@�*����mm�wK��Q���jk�oU���{�7��?���U�D�%v2="�G{Tq�=���`?qy:yr�7}5-��T���U��@Ӗ�|�Y-���h,�r-�{ۓ���\t
b¦D��7|Kΐ��)ȹ��Rť��C����T~x��{�m���d����;4ϻ�� ;m����f�l�zf�����?;|%L��\�VD����i[�h Qm��L��O	)���3t��E��=@�}����`XW�F��r�;�ҟ�����.n��K?���
ho�\	���������ȁ�&�M$���gd$!��)�}�r�()�ɼj�&�j���[3CPܒ�}!;z%Ԕ��ԉH��ܙ���� ����G����l�լkv���o ��e�N$��1T��`��Lj��PU0<訔�t���d{����c
	6H�I���X�P>���"W<#*�`���چG�p++2YN��������֫j��Eʼ�|\���aF�p%�+���Q"�"X��DO�'�:]�S&�����3}��f�pE��u��fҿn�&�!p8d�� �"�J���E�+�y���}&r����Xx�1�;%�)<ՈĘ��t6O1���g /���S�r[�Fh����<9��?#���9�"�H>cZ�j��WT�HXF���8�2��%[A-��(�D>rV�<7B�6W���wgDb����+@8��K6P#p"4�VR,���=e'���:9Wy�Q蟟e�/JT����U/���P��5���,;�R��}|�#!W���QTw6ύJ�S�#�3 ��Z�GPD�����XP�v���I�k�F���ޅ4R���\e��1�U���z2��uB�7���lL�T��#{6ώ���R�c"�<�n�4��9�o��-"�$sjF	�"�0uo����.ԥO�X��;h��{,�r�%: ʭ|�1����������b���������e便��|3�n����Q:�s��q��,V����8U��%��.����-� �=TA��q؞a�H�+�Į{�s�"�Ǭ�<��|���I��mOL �g�Q���3�YSt���Q�x�<,���~2�Ӆ�PW.�{.�V�$��tz#%�%R��+���<�ĵ��"	�V:�_���Z��&p��,f������^��{��[�2sD���}(��fx�:CP�e�R���;�gD�:���?q&��q�-eR��BoW-���mO��1|=���ջ]-��'@�R���p14���H3@-a�������#�lȤ��e�WZ%�R���:{�o�;�V�� �=��t�!���q���.��Q]��kA��ò���*���7ew���]��ࢇ^���Q1�V�"��Fh/H;i�-�W�&�/�fMr��1>�k�h�Yk��NX��TNV��:��X�NH��>�OB�碼[O����QHd��Z�ڃ�Y�)�$����q	7�K̆܅��"@f�������6dVZ��R9U��c�*_��50O�EΠ���KC[Uj��5C@�Y*H��a�M��l�́�s��<ԌTV �y�v��7�݁:�>�5T���oL���Y���z�Q�7V 6*ң�S�����r�>�&E�l�  ���4���G�ۮ��,���)H���Z;D3��O�N\Vo��?�&&�Y�<%]6	�k�ll{$�<�)�Kz����>	2�S���1d���V���F�4��K���X;lA^�=�!	�9Zny�h(~����0qĝ����u�M��rX�� �94A�h�������IR�6B�*D���됕r�����pYٰ��mI<ོ�U�ڼf�QO^�RF�Q=2	I�x��[a�衷�,[�k��j1}@(ovTr��IRA�o)+}�!YX���ГX�;�������Y��H�9D_�"�Is߉�x��Mme��(��~��#q�نw��XTs�uT��s��g�q��3�����9	7^�����5d�)�|a����f�fO�$3>1fёL�*��CA�Õr#D1/�y������V��:�C`�+���H!������;]xQ�/�~����'���/�[/+�%4�I��8���ۜ6n�,�/��&����������8����0S��� X�ޚe?3�
�v��\���nj�T�B��ez�cR�dڒE�,�ԧ�a��g�M'��>���ɃcH�Q*A��Q�{���r�uh�U�Ch͡�,Uq�/������C���l��7:3�}��� ���:���'	mч~��d�	�j!g��h�Y����5}ͤ;�1Q� �A*���M~��Tnu��r �OU�m�E,?�_!y�1�*�[�����l��q�n>�����@��Ȥ���9j