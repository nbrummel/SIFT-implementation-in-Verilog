XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������\ d8Or���D�q�}��>w�;%]�:����T(�% 
IT� k��͆��|�o4{	��/���EA��r�)"��n4�C��\Q2Y9��E�eK����y��f�݈pG�}=VA��A����U�ـ��Ό�@��'��0����*�a�%TW1K)䚱��d÷����n �w5��e�U:��x��i>�y����F$��c��H��qi�n��=94�/�fml\aF�d�a�f̶sE�n�/�#c6��h�WLG �M�PJ}�[�P�Gk�g��mT��/��A���>��~�&�Ȭ�v4���ku����g}mô�>w G�{����C!�/%&Z�������{\�%E�'����i��2�J܆Jq����w�n
���=��)_v 	fm۴B_���7)m���z����7v�]k�mby�:m�)rҳx�{��y�_}��t"�a��n�o���U��h������DFo뷽�B֗_��GA�}XS x��iw-�W�tVą���ú=�3�2�5�#f�j�<<���@�v|�Ʋ+ 0 ��I8R�z�d<Y;x�˭1�E�w�L�c���e�|�=���>��&�`:��S"+�m��p�F%�^�^����lyN��7k)$p�$�N���9�SB�s>�$��/�mp<
����e_]��86�,�����h���+^��6o+`������Fdcأ�����!���r�?�lx�vV'�܃,��V�]�:�ź�
ג��SHA�b����/�X�XlxVHYEB    761e    1770@���_��.��·O��J��J�[<��a���G+�R�I=c����B܎]<K�p,��S����̜RM(��������@�\PI���f{B��[���A?Xri���:���HFm���	���yj���Z��}��)������W�Sz��u{�^�TWm�I�H�E|��+�XN�P�b���i���ڎM��.�������Ħ����AZ�+a�ǳ9KB��:0ʐzI��!C�U̙"���o��yv8Y{��c�U́Ϟ���V&�l�+�(F����N��()��!Jk����A�̠#�ϡեDRS=(:ԭ���>?��'�`���:���$��v�e���:\�+ǌO�QѲ5�i|���x���>��F-ˀ�	5߷�>yL�tً�(��9�hm,]�B6ܔ猚Z�V�D݄"�6Ho|>�C��;�qL�n�H:�u�Y�Y̤��B�t@P��PlfT���7�/���H�-'�e�]�\@������c�6w4|VϚ�v�k R9:�+\Ye��5�J��b:��H�lw���7��a���eU\���Z�"YZ�5͔�
L���[p@���2�0��dvt�~D�����-fxN4��=���z
�̃[��*���K���vE�NV07	?���9/^�أ��ӽxj��{��vܡ�����	��L@Rח�@8�^�=�W
�
p�튿H��h����޿R��r�4?I2��%S�jtO��52�C��6�DC��POA-D�)*�����Oy�`q�%��W�k���ät*6���%s�3�+���,�W���&d���4XV'�Mjƚu�~ �G�g��#��ԏ�wFrm6<C��0��ąF�#(T�3��-R��·��7e=��.U!�;�z.0�ї����׉Om���2���]�K�t��:�M��	N���l٩�7�e��b�Ǒ�K�18�W�e�8< �橚Z���M��?p{���*OR�=:��ໜ��LZ/V�@�D�[��A��9���E��ݽـ3Qut���-�KӍ丌Dy��نu�!�1;�q{��W���������}���R�rWX��1f�^d� �6<c8G	ˌ]$�ćgl���uVﷳI	��FL��R ATY �3Щ)�d���Y�9%���S��َ���g��4v,���./]jxs��u��ÅF|�l2.|e�y��K\j��b�4��ۅ+]}bC�	6��QfF_��[�
�_��Һ?��V2�`�:3��3HZQn_��lA^�!��W� #�#��s�A��Zq�1?���A�#��Ik���c��ۮ1=��&u>�$;�pKV�����s��c�� ,�1ծ%ᗒ��(�)��:�j�mY�2��ҵ$\H������Hy!h��;�u��Au��-�$���PqN	��]�r{%,^CKso� QQ2�Rpt(�\��ty-fzMb!s�.�����y�!�(��&�&�=5Zwk�t�
Hz9���LJf� $KV�V������l���?������<�'=@zad�d�q��'p{�J��|��qtYipI��Қo���� ��c��.�h��	�F�UiΜ�ys|����0��;�2��U��J��fl��Vz������,_8n~��0���θ$�;���8���?����i�X|ij���vQQ�Ȓ����|�rݠQA�9f����U���{>a���$���9��;ײ?�XJoD�@fF�c�E[X~�!7���}l�moZ�pU['��:}h�iBX^����t�x^��Z�(�S{� �^���uK�{�<�&q�Q>�AF�-�^��CN��Zځ��hS&}�jx������Xk6�6��e�;zĴ1�An&��Ͼ �����؏���y�\���� Ű�,$�!�.�]lި�$��DZ=D
`��m��v�H��S#�5����,H�3+��/U�wr��)i%���#٨wj�ʙy�X��!A��^f�a6CV	/�kP�O>�J�W�yB,�"xo)d)h'|�g�����5i�+�4-�#���+R�3���S�I7>� w4�Y����4Y�����_�'$�JVÆ�mLd܋ L��;�e�����-����Y��H�݂�(�Z	���O�����f�R�b�ͥ���+�l0hq�1b�5"�+�Q"P4�"�(��i����o� �aAK��0�K:��j�C#�{}�$�dvvX/�p�D�fB����l-ڪ���t���6�_��]���I<�q�������f��r�_�q�m�-t�� �ty=I�̊iiQ�P�iv];�2?}�(�I
��Ht�&������#D���_�?h�%)�	���ۤ�q?�D���7;�,[α��T%��1*̆�	� �}LW)���@5ݙ�%�g���TopHZ��D�0>�����xՍ �R���"bU�<�D�"`a%��'X�)�⫌tgg�2��F�Kan�Quov�=e���	��V�z�J����������*�;���(3��k���	9Z:���e��� 
����yh���0Ij��?i{��ﻹ�Ī�i��:��S)�y��9���'`�Y.�*0���?���n��&�M)�)R�D>Cx��ۣ� ��~xHl��oU��ԩ 'Q^7�
ͼd)�b��֛妀��
 tU�J�<u�=�x��&ѻQ�n�D���j�#�s"Nƪ��d�z��>`��vL�b�[^x�����\�g���m
m��^�u ��J����e{��J!�sg|��no�Ia�V�nFk�u�V���ߦa��_R��#8Ql˦�k�&i �k�J�&���՘�rI��:�M��4	Ů�V�Jc/�����K�F"�	�L���v�~V�h��lJ�M~wi��L=�'��t�A�ǝ_	�8���l\��b��k��<��O��Ù��$o_M��������eȆ?���t���Q	�d�W�8��^{�^d|���g�#E�
�Šy���zU:$EP�dB�#/�ߕ�"Պ8�X�ݛ�\�4`i��9��s�fd��X�C�vb�pEl��~��&�ن����7o�l�!���C��`�|��&2'Dx���$�_�RBA���T �z�X���_�K���zޡG.ǳ5̤`
 t� w�фv%���NPy�({I"���İU����/=��K����V�71���O����c�.mN���z��7!�ۀVD�W��kg
�f&q���V[��k�\�L�aY 9�7z���<O���k�nQ�O���r
��w_i�J�4r(��*�^�U�Ҙ�3����c��B�p3���*c
L<P�鏿�׆��䆍�L �0�����r�wh��.k�*K��`������<%#!0d�,���#n9%�_���Og�<��.��_%�_�n���c���A�����}���@+�U#nySv�����jXw-G�b�%GUU�N>�+�5n����Ņ�H�Vg��K�@4�O���rvgo9*i2��!�F��h��7eoVOx����E:Q�
T@G#�#��Yq#�tNT��!y'��my#܌?�ã��q����e�H�D�wu��(AK�rϝ�Z���U��>�laZ;��r֥��΅��B��n�����ts�U��l}���2."I�3��p����!�P������>:��V:��:���:����2�i���S��Nq��Z�v��TJ�$�Ҧ<ϒ�J�1�>Ta��n�@�"��R7�u����xϡ��h�l�T>�r�Vm��X�f}p�R	!�X���c�"�Y�![r�C�� :��UIX]�Fۭ�Ũ�ËD�>�R��ld8~�C�J{
2�n�#�L�DZB\�"��UJ�)�������f=}�}����� |]P�o9c�ʤ��/[qXNH�9"x�6���V��]�ˎ�_NP�nA��h�Z%<�T4��`H��t�Q�Jt񐗥�2`��� �v�%k���n��M��w� O����Y����;Vˊ�2/z�x���P�-��zO��5��<= �UsX�O��I��$@����i.*��;kEs�զ.�o�s<�S٢P�U5�#���7��)��G��'-h`�����W�ͳ��+K\8L���w����؋�X�-�C����S��^͗1�L��DO�T0ʫ���.5�Q�_�oB�B{��)���/b?�wy���A(�~B]�14O�1��i�u�M�- �d���a]L޽%[{(������!�mD�4��R�[-�B���b�n�O�Y�� '�������פtC
��q{[��N.K	����[�����Xl��Ǥ�<��Kx�>���N ��o��7c�Z�y4��GA��^'������y*�tƋp���:�B��&�?��S�r��@��N�n^�����VnO��%7��1��s����`T�8���O�Y�n�+L�p��ꂮX���`�!vbGN��y�O!][+�]�_�^)_៞liU����v��I&�;�r�YK�9���^��[4�D���^:C?~7���k�����v��|2\���H5���~�b�{���Mt��Ddw�3�n�M�N����t1�A �Y�������"�'��Gh��!~�� ��T=׍�#���Qv���������v��Y{�:l2F�qP.�
�&}�w�������
R�K�: QX'�!_��;	M�6����=��M�W�wwqK��x2��P>iSǄY��F+x�	#�{���<ؐ	���U�X�.?͂����a�.-r�X�2����E���/���C��.�kH�3i����R�r<"����bwy��	��hE��-�ۓ
S1�38���(�17/�S;�����Y\��gA''U��^��Þgay��M��wy��I崻���7e%l�'�|.^��9�s�|(��a�L�X�G'��Ͽ�h�L��GP4�=�j)ڒ�c�j��}j�`|L/ќl[@�%#�"�����o�[�_�?Ȏ����X=0;t�A�T�sݼ�c;�ҹ�����
 I��!�m�|N���h A,v60T�� �KfD����Z�U�w�rj��_X��1�K��%};���ȣM}A4�������O���{�����j���O(��,@D&=H��0�k�n4�w���s���V-�Z¥#�7�����b6P�F�7��(`AתV�62��x��t\:O�c���3�˶�>y��uZK�<�RY���C�k����6�@g�U*�c�f]���Ǝ^c���sGk��k%��!�%r������J�.F��i�?�lx{���z�qз���6L�dT�e_;�l*�ԁ0X��4�т�?:�_?7���
N�X7��������紮��T�)�����4���fi���w�i]�f�|�紹0�!H����'������~'@p�.�P���~�59藿.���L 6ωUnR�(f����leS�(5lSpB�r��TsAxG�� 4=��q6��rM������k�z�t���$-�?�h���Mnk��7���Vc�����r���&(��K�*o6�+��Ŝ���G6���E�q�´(��O�xGm�U�(�4]B�v��Vq�g��y���}påZ�Du���*�]c�ebP�) G*i(ƪ8���CC���涗�f�y;)ְ�s����.�R� �eR���0X��uӮn��Ms�����P8 �q���6���g�z�5	D��草�[.x�ҡ,�}�-+tߐ�U������CW05��L��!��[j�C�����6kB�85,S��p_{��9(f��Y;��3�sB��!-��tc�2r��?�dko���x�ʸ����� l�XĶ�W�x��.^�����ױUK��t��p�\`���tƙ�+�N�*�[�jym�