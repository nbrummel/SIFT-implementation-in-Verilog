XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������#bX����i��^���G�U����'��1�󂦓���:!�{�����>��B��v�(U݅ �T  �����Q0�1ؒR�Əc�?خ��LPh�ӹ�2ÚH�ipl������2#"P���`o��F���܋q��v?��ڈ��������قRcv�8�ڷM�]��(0�qbL���]� ���b�i���S\��]%���s�+E�*7M���#�7��9~�OR�N���4���
j�`'�AMXG�]�r���v�+4�`��:��D���a��*�)t������n��`��J\�2Rh�i�(��eZ�@�g��n�~���,;-4 M�OI�Z���#�Qȱf.��V��2s�FB@�`=X馜�+ȶaul���I]Cd���5�W
��#�>@d��u�P��"PC���?Ovn�����3G�(�[-�?&��W�l�A�K���TJ�i����� @���@��V7����4>���S i��hŲ�n���r^�hih<��c����#�M]؉�U!�pE��٣1�K�'�-��E�,H�L��a#0�tP�����Hr��0���+�r�z�6�@߇�����JK��{b��������γ�L��*hD�8��o�f�,%����4��SM�O���A�-Ysdi�'9P�H�-���5��/	Z'?�‑���ߢF�*�=�?˲�:����׼zl�&��;vD����u��XlxVHYEB    5909    1550�ϡп�Y�?���2k�a��L�(k��1�G)�j�]E�W8YȝHT9�X�`�D�Ի��(���E��Y�$�<����Kn`��a#�����ܶ��rZ����(﷏U͏l6���v�~N7#2�Z�7�N��i�]�ؚ�Dft����O�� R���nQ�ӍX���+�]� �֨� ,)�~Q���M�E�*
F*��pl�.����2�W��e*�b�������G��xE����h"_[��\��a�C�%َ�h=1�,��~��{���ʘտ��s��(��
�,g\���fx:_aBBq����#�97��B�j��m�*��r� �@�"�ԋQD&#L�-ִf�2J�G�c7��Oz�4I�ɟ�m��p��싸�
�V�P�\�ü�WJuoƫ�G�����<v���Zd�/��̻���9�	mE[?���#ŭQa�L�H�Uլ=;l�H?�LMA��$�֜���$T�|$����4����ø"��f�jd�_E�����JM���#�ͯ��o�C�`��^�g�o���p�3���'s����r�)���,�Bt2�4��~>����'�eZyՍ�#(a�!~���j��+ �`<�����H[E$፨V� r��]���[Ş�l���dx���V����ʖ�TU���D&��)���t��"W���f��\�4o���mlڕ=�����yF�����I������l֌'����7���U*��݊�XCOw��ZM2�Ԃ���}_g5un:�y<��ӽ��퐂a����܀��b�oᰌM����R��Eգ[ǜ�qL�:/��Qe'�y�1L��L�m����v��g�y��T����)>Ag���w��m2L!��1|uO�i�u�Zn"N��	R�\I*Y�ɞr5^��N-�[�D����z��������P�C(t�d!�� �>��~b�������m���2��Ys����� �e�|�u��ڻ��V�W#c#���JD��r�o���m�0K�'��1Ҋ��+o�$���S��SE5 �dE���W+ʁt ���s"D�sD?O���K;0#�}�B����Ad9��Y�Z�����:�[�v�0w��$�� 	����%оG���ѹ�c�������9�}谞��������_^]d:
n���&����X���o	�����W�X�C����羌�u��Go�[7y��,1��`�cm~շ��gNG�a$Cs'U{�ikͣ�������n�J��y��� I�/��e�Bl�cH�u������@¾׃��ő�2���Or_Cs����$���~�MF|��2fi���Qi����Q��Q��@���P���E���β���A�.1_Jp~�
 JصV�X��sX��/%)@��e��nl�����{O`m���w.�j]�s�H=z��6EN�qC�H_R�Ww<�����B�b9Sk�'��k���Ə�E)KLA���Q �U�3�j�b��YgW�	-�����dmܔ����0{�����u��<u����[He�Ybk̶��o�x���#��	浭��'t�W�Y�e��1Ny*�旾S��l�ٿ�ɩ-W��E�4�R���>�� �+��е��<���q���5MF�O��tn�Ebe��z�?fx�U�*Ȧ)���D�h-�bd&�=�s ����B$@��L���ji�Bt�M$�lɭar�c��o��eh����~�����M�%��{��F��6�J`e���?oFZ\��u�n��G�$�l�=ܠ4>aU��E��	TZ��
�ߺ�M
�S�-y؂#K!n�ͽ5�s2��l!�c�{�N汭����k�P3�d���xp��w��I�4��\( ��4o&\z�!�5:j��(�		��.��~4Ҽ]��iv�H}#urj�KBD�1�/�uA���yw��~c&��^P�5���G��AA�f�� *0b$��U8X����flm�����~0.�(�Z	�j(J�*&�3��lj�����:^lN*A�<���%�J����W~���f�� j�� ���;���uO蛣�u۪��#�|�j.͝� �MNxE(A� �_�:&`�
b��B�A����KIx eSOt��:%����� ���	��.;�猛���p�k�An�6Sq�D�n_� QĒ�Td,5���%�Rv$�Rb�}
:qG�i�`��1G�Hb��G�vɑ��|�#!�C�b��a�o�<9�V��DId�
J ��@g��!��6fL��7�T�=��YM`Gt�el�Vӷ=�A|�Ǣ��UԌ�\?�a�C�lko�Mu���1�f��+��������k�/Jޫg������9�ix!w��kb�p'(�K	]�a�gU�T������3I��'sAd��
�%	)i�&��K��-}8g�:�u��V��4y1b�=nF��]�i�<�S	7�u�( ęס?1���*};�ʱ\*�T�1RZ�+#I����<۾�b�KcR�]����H�$�S���:��h�e��S�/M����!��^��C�����6��'�%����:�`�"�G��n���A���l����H$�'��M ���#��=�"�A��߫�3}�+��.�D�y/�\T�E����S~01H�=�"4_|�+37���	>�P�$���]�>���}8�-Jb8��[w�d�,R܍�od�^�n����,|�z�	��\�����o<y�;�����tE�Lyf�F�7ԬQ^�|o�J:��K���ҭKH�ȖϹ��@R�7N|d������MIUoKy���2�	�z��7�´��֋]1"+�W�)s�^ۄl���WPi6�x�p�=b�nWza"�zr��IG�ܜU�A7`�k��R��bS�(t{X8��B��y�v·�iI6l�SK����J��T0�j]vH��#T!�@��A�_�.X!�j��5^�?Z���Z<М�iwA����a��46���#Da�5�v[�q�Cr�Jn��9=\Y?��"���=�3j�4�����!x��ĵ�1(K�pf�)��o���u��O1���j(E��E�E�Pfr�վ2l��2�}�e���iG2���q~��4�h��J� gq�b�n+�Õ.����q<�{Oz)h�')�E��sTz�Qʣi���zکT�n°$FE�qS8�S�ͽ�� x��Y/7NA�n�����'7�߱D=����G�a��c��ڎ��?�0��� L���0�:x�.\� =���y��&�ؙ?7��!���z'MG��M�~��h�#�����$��_m� a�p�tt��z�$RΞ��e�t�e筒2�
ډ�fL��Q���mdn��j��b�.A�q.��n�s�ϹY�>�ިB_�l�ĭ}_���>��7�9�Q�մx==V�<2?�V�c�6�Uq覫ߏG��J�DS����K�
��G�n٦�t�jQ��4deMH�*�eO}���~54��ֶ	�,���Ɩ��F���J����ֲѩ �g Ă�K�1-"��kq��a�[�~}��?,z�)��~�I�k� �}�=+�R�p8����uT*��/�1n�	y�i8Df�v�4�Ҝw�l=�1U#�]t O�����Go������^)�c�Dw�w��J�i(%�۶&j���F��'�x���� �"�������9w��e?p��L��5)?(���Ʈ�@X�s� >H��bU�W���E��
a���xG�at�VY�H{���2�"����$8#�PZ���{�N���G3����6�쯴��X�a�y-_�C���@ss���y�?�d�ن���L�݅u�����GU��Sɘu�CJ�cZ��O��fs�3��W�s�Y��n���o�k����a=�M���D�2<L�)D�e���n�`{�^W�^�~AQ:�
v�)4Қ�n-аI�����i=ƆH|U�0� W$!�m�K�)���j��¤-�o[#{4�<g�g��"g�n-}"02�g�A��F�i�'��l���3�Jrx���l��I�I��H��Y��`�/i����@�Yqf]z���;�t�u,����yLˣ��*�!6�O�41is1�eb�%��r��c�p�:�ṫ�S՚�.fQ��X��v��R�גKQ6��+�}�?@��C�j��S� �៳Q�],Iid�;�<���&�� q:M�GVX��+�l�*�n���dԛA�39\�!�uW��u�������3�.˞g��
ј5�!	�n$iF
]H��cDz&�˪�j��R�c�`߷Ƅ=kʫ� =�΁B�,E<�|�&����<q~t�Y�;��ܙk�]�d�f���� Ld����I����+2.�	IuE��Դ�o�����X�˞�/N{��?P��F�7*ґ�.xj�.}
�kn���L��oZ�nZ?k�}A�״�^ߚޱ����6�	w�ޠtۍ�.\�&��>U�|������A}�q1�(+2<�S��X����E�i〽��Bo���b��R��F�q+��Qp,��[��m��n���$��@cq�L�6?����u��e(�X�r��٨Ç�	6��_�b�a�����x�n��l�VP����S��y��v�!x|���vϱ:��X6�h��3u�策�a�O}v&f>�b~��V���߅l��k`�̯s���]� =��!<�	��bM�6�A�ƳJ3� �΢�c�3$	�3�	:���_a6G������b8�ې�>�U�������#�<�����1v�l(,�o'X���P��o�,v긮m#�4�o��-�r��⫍��:XBS����p3-?�ރy��)IK-Bfέ��"���J��x�ԋ�������|n0����.����5|@��� �U+����EA�_3< ���Lj��F�Z������1qۥ�������iP�ݨ��A����	�-I�Ƽ���=���`D(��#��+�E�v�u���[C��	t���8 �0��d�ڦ_��e���<ߋ�t_~K֜O�n��u�c�?���'2~đ&М���7�ZA8G<Z;n��r�_��u������X���I��t~���|��L#���&?�}�l��"��NN &���Ho��Rބn.v��xɓ\�i�<[V�7J?
�����+"�4�)��Ewا��Z�@�  @���N�M�)�z�z��x��^G+��	t�Z��>6�Ђ/�G����+%
��M���&�O;SsC��,B��I8�|�,�U��c��x$� ��N���,�����ҏ6WE��<�� �Z�I��g�~��������^��\	ǜ�tΕ�#)W_;_��0B֔�3,