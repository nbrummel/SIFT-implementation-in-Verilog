XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-JZ�M?M��._�'���5,�I��O�d�y3X*5�-<(��O��{�vdC�(��Q!Jz������.D�E�p�VK2"\�d))9�޳�(�s��_z���k�H#9�9L�TdV2#���;�W����C.��[��k�mu��c�&J��|�*�fI�Abl�pa킀͜'4����BD@��z��Ld1��#<�7D���!Ckyf�bU�)M> �y�u1�^$��M{��`!=n� ($�P��8�3[;<
�0/��F<���G�w{n�ۢ{h��"�� )d�+Vj���3W�i�[!b��IN�]��2LF�O���?ݐ��%���(�o)�	��+�� ���Sɔ=�U�ˢ_�j��Ā	�����XU�;*�w��xR����V��P��BJ=���D�*	4�a����Yr[�~,H(jyXKg"��I�ߪ������p���Bz^)ݸ���yٚ��4�a_�ӷ��J����{o�|7��\�3}|������Zo��.<6��'����0B�s.#(�DebI
�:,��/6C� �@�0����,[>,B�o=��+D�wYw�}�G��������+< �:D��|�>�/�iM����\�������3�C=��8A�u���1��_���I�7����������F���?��99WYV�9�y���hAeԆm��k��Y:VE<����5�c8��ۯ���1��z%V�ֱ�6���=J�eo#Kf��XlxVHYEB    7744    1780
�E�ʭ�K	������/!�EeU�'�r���G�y�e�R��4�m������m��D��R��|�Cԝ��-ܘ�G�s�!�*X�����#`���������_��~�8�rq�b{,O��3�7�ׂf�=�~X��3ځ�M`����G���{4T�-Z=
D�<,"�m���0��L����]Z�9g`���Y�J���,���3�<�gU�4Pe����d(���b6_Q�MݙI)���n�Z?�ʪ ��*B?'�@������4����S�_��(!���#�������1wi���ʹ��*��K�q��}�aAfB$��SI$m�.������_�KY��5�3�o1g��ŧ�%���`���;�c	-�� N��?�f�[^p��hԟ�e��ɠ�bH]z���Ӡ�M*8�m8
�i�?N��Bx�b)W��9��X#(�b�z���A:1�
G�0!���	�03X����%ȼ�2ܟ7q/T�i�")�e�k��;n7�d��R��=��K"����W�w�K\�3��8.�s"i��K�~��,[�����bm�]� -��B���1��$�%��4,`��X4G�e�,���c�����Glyz8�2���8��2`�ʎ̄�� �i�I���HK��圇��ʩ�>`u ���ymz�7���g��ɷ�>h�"�#�ތdѪ�b$q�Ӝ�sJk8X�G'\R�Q0Ғ��S���i�?�
x%-IyJJ�M���`��>���E-�bE1�$���I	�ǀ�����l:g'�V���9���SI�K̀�cN�	+�wx�����%�P`���hDI5���p�	�ͨڏsN^��؞�@A}��䕣�F{:K}4��h�{�����Ypq_G�`���F0��,�-��{�9ǣ��]�	�n�8Z�1�ݛ��4(.@lɲ�l��;ْ��F N(@��2��$;_JsCyh��"���LU30��+�ǟ1țȔ���9u[��=/9I���+p?����"��Z��YުU�a���&I6�ΨmͥW?���O���o�j�l q���ڝ|�������a4.#����{.���\W�+]�����bq�¢c-S'�;V���ɐ��X��(�4��w����B�i�mX.ۼ��6)�A}3y!¸t�X	Pe!~+���o�o�Ţ|�?i$�M]��f��i	��@ao��}���3k��KȾJX���8�4��'�ẎGĭ;^��]�_Dm|�d0���^P~��́wW��X��o���(�t�'Cv[@o[0�Z4�"���d_x5���g����ԉ˜�sߣOt�=���W)��>�c�A��rGxGԋ�h�S���dz��^��Y��%!�;�9�x��d���B�#�K)�.�W���w���5��ֲ�i�f�`(�
�1�T�Ӷ&P�3$�k�0����c�3�uι�V����_{==���MJ�m�*���͞�Q�g3�چ�PU=�4��x[���Y��f�0�&����R�Ce�@�����sA<���Kp	L����S�7��2�?�	��7gK����x�� M1��ѫA���5���X��E�30_�����L5)4v��4�$aİ�ۙ�á]�j�u��ҷQ��¨n��k��l�+1{��0��)�+3�k�)}�
���<ާ�U�����@��Z���]l�8+e���L�얜u��ĩW�<�/�=�f<����/�y�hQ�VҖ���R1	��]���5>%r�������![Osa��\�7���S��/_~��x��~:!�|���]��F�ރr�u�Ϗ:�:�t�s)���I�bA�7U8(%7�����s�U�͵J8/�Mi��k$���Qd�]���0����Zxwk�B'�2��� *{�l�B�D�-�ă�9��}ң�Ǟ�w����5�H���u�� ��s����{�"nuQݼ[n��Z9�����8��������'�G�	��;��C��t;x�i8����v1�滆�
.X,U��n�Qg�~v��>\`x�̺��L�����bI��:<h���ZݕEU1k2vP�V�k�d�<ˬ�9����,��@E�XU=�8�v#���gu�Q�jV�B�jRnr�N�8 ��K�l��L��� ��ʫW�뗽+}Ձcϸ*�x�����z#��^qW읁B�ɺ��O7��H䎽h-ݠz�Y�D�����K^�:"�����%�s{��A������������e� 8s�<�2㆜�A@ 7�5��� ?e��� �TC�L�6x��߱�YЪ������~��Nv��8�1A�!N.9i
%\���΃H9\7#���X_'��!4{~��^5/����g�*�ڡ�WЂ��,���~ɤj��|�:��-���d,��
20�<���U�E��rl.��%I��_�,�����S�5%$˽��L���kioi]3���љZ�����b}d�+o�tIq�F�7�s	b��^N�f�EB��D�vþ�c1A���x�O%�J~AQ����Ц����NK���|[c�}f�M�g|�Q'�]WnD����$�D�:�О�~���`�&�$�5?;�
����Ǆ�0��Q&�jr��H�?j�-V�|.MSВ�D
H
��z�(R���$�.ڍju��vc��4��2�?G�/� ��lj��J0),�-ܕ��4�%��_��O�6�c�x<�%hU�]=Bkr�\�[�}^���]�#��
�j�>�ԧ�P�(uL�gu�}���)I���꾏��	5nSs$� ���kь �#�7���h�Îd�ʬ���� Cn��fڹ�����|d=�S �چEo��r���\���`湋u�k>_ÿ�bo���u�Yڻ���/��A-�3���@{�1��X��ɗޔoO���<�9ȅ�U��1&%�=B}�iI�;��5�f77k�O��5��$�U��᠂��84��{4�2���l\=,x�6w���|�o-�'M*�]p�vfZx���q`L�7��wލ�K�|i�IQ������oΰ�����t��A�SK�v�����(:��W�Hځ��}0nT�I��-f8Zd�[�ؤ���O^��d�.�������9��a -�&���c�����(Y��od!Є������§������I�5�k!�ݿ7��,�^��]g����3S�v}��g&\�i�{,#�T��2J
��wU~#@�3b��<�uQ7��:o�Ki�7]����4F�˳�5<mH�I��F��џObT�-�2�$,J�Ȗа�hb�w��D/��{SΩ]�EF͉�;|�b��b�������ޑR����&+�=L�����Y�&�6!�Κ�z6�u��7�2D�1�C���\�O/:�еoM�ʝE���ٰv��:ũ>%��/l���6������n�W^��R#�J��(=U�l���I-��jk�z���r�#�������k����>��5wr�< �	U�0B�R����>��4�f Ù����Pu�PG[����an+�hB
�[؜e�%Kj޷���ϧ��xpV��i���7����G� �aI�1��`��H|�x�&:��1q�,K���Nz�ye Xyw�D)UL�lᆝԛ�W�XA�޾VV8��u�f}�
On��r�P��a�
�CtQ��7,HxϬ��mH��u$��.���/9���X;.���F�����}��x��dA������Y�_�;+����蟘Ӛ����X:T�)��w�=P��s��Yc�}�:#.�.[3�����h�lA�����adB�P6?k�kk:\�^���Ĝ�1kB"�_�W�q�������������"�������Z��6^�{�	��X����p��W�ihӜM�5�sϚ-�F���(Rr��6Y�r���},�@�.����,L�2+�N�(�x�ld+Ù�
wR���n;[,�)ʽG2��0�M;_�̇���˔�u�y�])���>�����r�j{��ZT�pϖ&���ls܌�3��
P�����%���M
��~�a{e+�L��`f��-��}��O�B�	
����Ќ=M���������z�eQ�)�_��-l۹}�k��2 ��=�~�5����iDږUQ����t�����S�i�����'�mm<8p$g7��y��t�!pyq�QS��/�.ǗV^r!�?�m�3F]��8��ҘO搸,�X#r>σ���
�DH��S�39��1P	!Q�fS��	�eA��3s-���I����ऱP��ժ4Y�'�~pO��4,�˖ё�!����&1��FG�1kk��/̼/�3�؄��'kVC���8�:�l��PO�i��o�X#V�r��Q��:RC\��#��r��q�Ȍ-�6%�2��e��9�T����m ���W�u��(&�u�0�řآ�'���;r��O.Q�k��^qs�.M��e$┞��m�js�ٽE��w�~2��~R�m�J�G��i�;��y���h�V������<��j�ǿ�V�d!b�D�ԑ����>��uCE:���ɚ�ӯ"��(T�$��lS�21�8����jL ^+�U��x[��^�V�9���|b��ޘ���3Kf�;�5�j댴":�ԚH���udt_|�G�6Ӏe���$�Q롰1������u��e�l���`Lӭ�+��$�"K���l?Y�a��j�"h��).�.t��$�kI�d��������=x�ze�8�n�p�،�e~jYS2�kI��[9���k�W�b����Û%ڔ�*e�n!g���La�[31ۇ�o�\�I�h�	�)�aO����>����m�\��Z`2@=W���5mXj�bcV�w�Ύe�����t�������[�p�a����fMs�՚�fy�8\�p/�pm�RE��������^��e�n����]'>�����8�4�2Ӥ�h��j�S+բKu�v�
Ƚ֧�bF>2�ȵ��}�Z+��LL��������w�J�,�شt��?�z�w�#�^�D�@% Oke��=XI���5$� 	�f��ԫr������|�Ǒ,��\����I1f�%q��2pJ*,�E����<��Q�n���i	���8�O��h�Y�A�'��l�S�E�����%I�
�Cs�p{6� ��<	'��ߐn>�(a�@h�O=A�Q��K3�>\H�{����4��0<�\��m��?u���Q��u'D#���c��ȿ��si����}������r\@궒7�'}��s�B܆�Yt��$.���s��?<H�Z�����f�n�C�ɂ�մb�M�(	uVb-~S���)A�� �>��� q_��C�"D$)"e�[��n�o0״�A��n��ǺTY��+[�̆�E�CQ3Q
�+r�p���'<WM試�������OI���_��C����'�k"�X��C�I%]͚��e�����(��	�**�}���p�\�RR�T�(�<I�=W�gSw���~����q����9ɱ/���q��@����zҧ��n���p�a��i2���%��E g��W�Z1�x��[�n�5Ln�?S�{��������u���@�n�6���˭�����R���QM(޸�h�J� ��*Y*��4vRl5�h��7�J���jt�X�4����
��҅&����Sn_$���&)B�f��tk�x������ST�Eem�nѥ�V쁚|��������A�� �E��\s� Be\�u�S���xy>�	V�R�k��i3�l@D�S�\Bg��<�uf2c@"S�Z}=�_�C���t�S9y���-���WTcpŸ�в�$w��e�Q�Eˀ�|�z)h�?|z�[���V�Z�x_����}Oga~�c�8㨪.BT&�QG>�*߱���?�Plŷ��ެ�