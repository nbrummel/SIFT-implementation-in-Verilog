XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x
qPfl� 1㌍m5���d��؊�[-�8a��=��C��o/�50h2�6�d���¯���o�w�O[��m]�-ed&�T�~X���srwzK3Ӧ�U�2�?���8^�����8";Fu����#O"��y�F�t�Gh:�P��q|�\̕���X-�X���F̏9��B��e��ڗ�k>��6�@!���RH�z���Au}�? t>�����H�+G	��� BoC��'���|�4'��)IA4����_�|{s#MQ��-fO? �J�Z9uq�T��@��T��@���!�T����7i�-$ �,�X���Z&����t�,�	s)2�e��ƒ`h}c�F��y{@kdiF�J�7�h��͙_��Q/�4������ˀp%���p�oK�
�J�B�I�~͝��Z�˟����_�U� n�3.�bh��Y�r���[����p�'�e�b5�ػI�"��B�lZf��4��`����/�����,+3�Г�D�?����K���|�}�+LX�&,��Z��E��ᘉ{������uoӰlOb�b���<,Ń���s{7�Ȍ�����M��R~�L���[��H!A(��q�y�?��$6"�Cq�y(�����^��=W��G�4��;Ҍ�"�ׁ,��Tp�pc��0�X��� U�K�����E#=UJ��rd����R~���}�8�=��䚽G|_���-ك뭓�p~��e�|#0�i�ɪ�i���U���;�A��XlxVHYEB    aa31    1e40*������0���	�n�3vS�^�i��[L$��h��L�F��Z�l����R	~������)ǮT�e�T�=�R�<�a�#���H� �y?�d��c082yT��ph�W�>	�|;Ȟ�Kg�F)"M�-;�(���$�NTU��W"v4w#�����v���} E���3�v�$*1�O��;��F��@��R�1&R�[&�}�C�s�`�Ћ���{m���Տ`�E�e�?�U����Q	#\�=�T.��4��Wn��|g��M�����I�I�f�o��c�P�����l�?�ĥ���Ỳ��d��R���sWM��Ѥ��䊌D�$B���X�xԖ��5�b�z�s޾�)V�c�%��/X�t�(�����qp)	����Rl/���� �cø_wK�R{s	�c�]��ti�t��'��4��
��t4y_�J��}.�JB^;*�c����=4mĝhx��M����UK����ls$'�6�F���l)�ԅ�9L`g�h�3�ġ���7�4Q��Q���~J^#KV$���=��\kb��X
�����>3'�z�}I�E�~��	]
��?)Uj��v�ce'8k�
���P���=O��Zz�"
J�35��Fȍ||��7�Ĉ�iSf�� $>��w6S��T~b��i�d������Jpeԋ�B��#�tZ��EC�ZT���A�&'�֟GGJ�%)w\�����G!fU�a��̐���8��\2�6z�D�ez(;.����U[Z�i�=4F��t]����n.u�#m
�����S���˰�W��&-bt��K�_��r�~jp�S�b� ���#��G]��2��GC�"Գ��U2"Z�r�"���m�T��������	�yڱ���R�gȮ��KU��O�6fSV�Uc�j�uRI��^-H�,mwBb^��zNBY���l~����
w�����u����x��)(a�kl&���P��fM�CQ� �e���,�;F�h��s:>
p�%���1��>ᯛi��*P�۵�n��SZM��e�����A`�V�Y��k���W��<�
w:��)1����8#�DuHJ>�I�I�"BX�21zC���X�� ��r��E��I�E�8S���?�&B���,U�-�*���F|�0z\��5��ŋ�S�?�Go��fk��j�7�rLO��QJ#�� �I��_b��,����E=M�Mʡ��IG�SIC4ѕy�%�h�)�~�I�Kv�0���Gy��זOPt�a4'�|���Mx�O���L%T'�s:������|N��Z�9p!�)= �cm�x�G�J�^�I��B��qO'+��+5��
O)Nv����*�`W��[�[ǖ��Ȍ�~x���J-ZvB?��D"�xS�FB*���M�u�i�!0�lAҽa�:������$)Z��Ϣ���N��'�_Xĳ���uVw� h'�`�������TIo�;� ��R�@�[ր���$�^Tf�rP��t������yX;d2��� ��9GNAqw�ꛗ4��9���	�6fOy�o~�m~aU�����]�sH��Nv��]��L���: ���ۓ](���|7\JU7�j�U����v�<�J��ИD�vN���Ԙ�sD������I�e$�����Z�	�����Ąiu3���m{$��P�r;�O�I���e�(�r�66���$v���6���ai�:�L-O�So�___kL�|�-�����+�P���@0�$���v~*9�WEz�E8��J�<��!��j��I�Oٓ�0�{1��\GZw��Oi�O�GjT[��.r�M�J�fU�w�'����<��79T�m�)h�-�+(�_}B�"��7��s�4�2[]-��q��Fc^�I^Ϛ���\���1���nkY.g�[�,��*M\k�s�~ۈ�r@�2����q����8��T0�G���Zf��5"q�H
�[��,k���@PD�I�p�Sr��sZ���X̀��F�:.���&{�S�񜽍�}ɕ�>/��e8ҩQ�G� E�eG�jbOo����ôS����\*�:'��i-�uq�(�_a�@������\�J�Wu�w���ϝ�;DPd��h;v��Q1���y�gLt�/ŻIQa����h���B��%�c�Ǌ|�~�)/��TD|��r�b�[~)���@jB��-���_"<�D.&eZ�xV���̫�o�^ozy����w�N���+����N���-�&>��|��R~�e�8*M%C�r�O�d͝���4^�FC~���
�j$��ߡo(�Ǌ&<T��C;��܋��-�|F��l� A����"̩u�j!o�pM� .a�ȗ���Y��D�G�SM Mq�I��GZo8.��J�h�Q�"�=��~���N?,����LxYg�<�U��$rvأ�F���5�p.�U_���Ѳh�ưx����"�{�����'WI��B�0ne��y�b��;�C�#\�ay�� ;CiI"1.���F�Sδ�Zp7��KH�&{�*T��y��
��V�}�׋4�ҵ�h��#e���{��Wn3�ӗEea��-WrX��OH�δ��6�S8�r7�
,�]Q��r#��2o"��~��1�"qc�w�]s�HbR��{��j�j�]u�i�kG�_���k���}�����.����V��1^�ro5v)nE`�0�-��DEO����*= ��Qa���Q��*�?����Aֽ�x�BlcИp9nO<�+���<.���'�N)I��،߰��W�=�|�.m#j*O�,@�Q'3�N��*,��R�j�=ōUB��p�v}�c�U�t-�n��6y|��6�z\�{d�u�ԍ�f�.���raA~r,���'�1��#�.B��16Nv��a�-'F�@|����}�|ƪ�T����^�hAA ��혤��'BL�!* � ���>/���/��+�$-�욳�Ή
���KS�F@4���6��e1�}�q�Q�r"���.X%�S���Y�K�C�^
s�\M?8������S�jIY��qܺ�l�,�,sRӲkL+@��d�qs|Xڔ蜃�%�Vh�(�;�a��>��rT�5�=��L��maTYMJ��t��W�<T?���sZw�Wt�O�FS|��J�;OdT���oc����zG�nʚ�D�7O�� �7B�,Z��ܴ-�:��Ļ����CD���3�\�Z���-��/h�C3�\y��
�[���6�̦Zt�}UZ
N�c�|b�Ũi/	*x�Xj^-N��p���"a⡘qT\��LD$Y�sX��z`�5�Ճ�D���3��Ч8��MW$蠮���E(��Kh\ʿxc���(�r�k�W��\bi�c�ڑ�^�9��3�2��������tj�$/�6�5 MU�m�?�-���k�C��:l]z���@7׍� s"� �i~�?�#89�-9ğ��&>5|[�%\�X70��EQ�����#��r�ȧ ���jw����� ��������ǘ��#Ձ�ѩt���C>s�F��u��;|��eɠ���s3�]?O1���L��u{�!���i� �Wq�j����!�,�:,o���K���ΕߤlvJ'D�"m�ܙ(`�y�fa3Hg����\nЭ��]k��hCDJh.U"�E�y&���F�4�a��K�$�������<��J�1i�V�Ke�(Vo�F����+��f��9�U�n�.P'��D��	b�`���8��Vo�?�d$�dJQ)��D�!@S�m�D����7v�~'�?�xĤ�y�;�},�R��V�m��^�i�"�M*Iz�\U$���gW/��6r�3�X�{u�����'&��O�~����o�ϡ��	�,r�{�WYi:E�J�Ji�"�AC���/���yy���F��"2���!�H/[�%�RW�w���,���H�=�:6����z/k��̆��Ν� H^���1g���O竛� ;����j���._�J։C1��'�j����ɚoaz�_��)� &𢸧��l��<�A�$Ax����Y=���Sᦪ����8K��{D\��$�g�#�X�o��ЖZ?�$��6�o��2���Ro�I=	�Q��y��Y��jrꦕ��J�/��V����Rz�i���g߯`��i�������;�A�:�����%��g�#��֖�u���Dqc��C]0�?���;�A�ACɀ��Z�������˧W }a?g�L7�����`��y.Q��ɭ�zW�j P;��4*e Nl��mA�;ą�l�|xA��5�A�ċ�ע�p��Q��e�|�^t�K�&,�^�Uzs
C�#� �c�n'�l��6���O���0�{P���|]Ck��$���y�י�`At�w�Z=l���O��Y���������w1%�� -}�(�щl��i6��kᨌ,˟��-��I�&�DC*̫���΄�� 9H��^K ��Z}�?7ߪ��u�JM����I���n�v�����7��z?Q�����Ķ�ŗ�NVy���	����G���R��B����Բ)��҈�k�,���f�h�4z�="���{�v��z�#�ј�i�=3&�ݽI�Yv�fC1<������3�t�̺�r�<ݵ���E���.���~�$o��T��dp٢��I��SC��~
���3kuJ ����E�w 9F)���r8�/Ȃ7�#�F=��?����$&�j4a�B6�cB:�O�~�����6��%��Go���>��7��{��]�ǐg��������"��%�r�-
�{I���Iq��0]eb	B)N_Up?����|r�k�{��+�
�bC5:�"Kb%ԑ;�k�C%�1��-��Up��kac����ՆO�@%K�S7]|�T��9���%��9��s4@X ƕ�܌���h�i��K�C���r �	����yIp}�B����N�
���c�*�/<)�E����یW����Sw�Ѐ��o8bx�`�ήOֺ���s�&�������ڮ��q����gP��h�V��ŕT?�o}?�7�MM`�"��q�6��K4���Ke�E�N<�(��x�jy�RP�| S��h{�&�y���.����jBj3�H ���?�H �.M�t��(��Wgh����+�vM'�Jn�P��Ȍ�
�>G8��@�qUU������>!���bACB���ۃ�<H{��	ם�{'�L��y(��o�-��=<��*�b�������eh.Vi�oʐDvI9�Mmg/f� Fv���N��O��g�Y�C�1�a��Jc� �4柆)�g�w+P�ܶ�Y1�)#��Nz�,B�
(����P�:���{���F(�L������É�$I �͖¿���ݩh^�<�W��A_qQ�Z�I�E�E�W��o_U���]�R�i�z<G-�Zl/]�I{�Q{�gߢ������˹d�`2܈��(�k+��A�ex���2���	`����1"��'W��5=�w�A�?0�8�k���_�@p��|�up[���ȭ�,ġ��7��b�VA{��ya؋��48��p���ڍ$��W�@;coF�}As��f�E�+)�:x��V�>zh@��<�΍>#w��ҷ<D_'�!?U ���{>�$�״J�*��8�f�k�`���z��
��B���d��\��{��kfP��bN�bq�';Ȑ���_���oxL�kK�)��1�/x�j�l���h�f��y2gت������	�g�&�㩩��� VT���~+�uC����D�a�}���ѕe�}Eԭ����k�:�f��Њ��hJ��c��PQoa��8_��siq����/���y�[?T��%H��M��'��BP00.S�5�-��˜��DVfS_&0h;�c�~��ewQagb�9+uqf�����;˒A [%e̥�����Sʆt}��A v��#J��c�@����.�p���L��M�ż.��Yx{j�#�_vB@R��o쨟 �?�Z5�@�\;����*M�v�FSч�La�d�U|�5��e:��.�V�}5O��M�(
/hՈ\�5�{�-�B�:!ߺ�*�V�c��Ӵ�F���2���E#R�mL���N��{�cd�$�.b��%=7��rr9/>�j�֠XI��T8%^��'³C{��(�����lL|��~�%�V��[?�t�7��N�Ju�2(�3;�3,+�0yI���L&������X��2��줽ABiʫ�Z "�~��_ҕ��4&�����f��c�մ������OI�M����s�[�J�%�c�c~6��;r͜Ғ}�1_���~���j���m�-3KH�.����>H��%��G^2�%o�����L�� qo*��h;M�$j�*.�o>�0�{F��f�;�>=�j�l�}�N����m:w����W5�5�3�"���z=�tɢ-���������Cg��.�S��!$���Γ�����br=�?��&f_~�
^i\r�2�Г�;4��|�6Xt��&�g��H�����'�S����b9]Ӏ���~��*ĔAzHT�~�\C -�ΝK�Ja-�j���N�� �iń~��'�D����|�⹻߼C��n� ��!0�u���z|�������r1Z�}�+s�̨��(4|1\-a���S���كl&��F�)K���e� ��/�����F��H�[��p${n�ǥ�Hκ�����ż�s�_ʹ�뀅ՇJ��
��䣠w�5��	|XgH�us�B/�Y���p����\��YC����`O�b��Q�&���o��@3���,�I���u g�A�����/�XO���'��x&��ጩ�"�u�E�Zu	��&���Bh>�u������tv�T���XR���Ye� ���乲�q�"o�tμ(�����L��>#kI�˳�;�]���K$��u��������N+�t�IR0�6Q�TZ\�	z&4�j�M��Yh�}\n�IĂ(�G��l����4����6���~-�8YU�� 11k��2W�u�X�s���P5�V���c��6ьn��.79ɏ�Ir �1'�7:�C��-�n���l�/gKg
E#nG��f�a��R�+Yد	�>*,�5zz�WvfW�KK+�M��HO0���l���Ll-����zRt�L�J}v̪�y:�?��_��1�lO�<n�������R���}�u���y˥�A���N�ӾI�m��n�(0qr�au�sz��_d���2�c��"Ш��ӊ�����S���(@��"���Nқ�:(���%h��Bu�,���.��_bη~k^�{�ĸb����U/�ASI��%��6v{n���噛�Y����}� ��-���v!��Q7z��.?� 2� ظ�J ��/ 0�?�����t�E��X�W��zM��~r ��c��х0z��Mg�']H��S��H8C[KNC���u~4��&%����k�0]*8@Vly�/��y�?��Y}^H�sC�^٢�ԲA{AZ(=�X�N���I�ʲS(�D|z�����'3#[�VAj�Ud���ޑ~�"s�E�m~