XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
���O'��,�U�5O>�C����M|�.�/}��惬����z�kү�m�ա�] �t�A2�����p2��M8���C¤|�w�
�|�D%�߷�Pe�#���)%4�J�-����ِ�2��)����Ś�F��
� ��f#^��`,�5��(��*!������7�����J��n!��'ɇ��!b@��=��@툼24�q��<ip�kl�m`{����yPn��I�]�mۃ�߅hS_H3����Lϱrc��:"1��QƧ"c��VYI�DWQ̚���P/��(�5b՟����$p����]wૅh����� +�]{���ԭ>�u�<�(t�!�m)La%`��Z�E���+�����>����SJ|C�!	^��k�Y�ጅ^k��:K�T����Bk�����x�k�j�X��i�@R�T��Dւ�ňDM�^J��(�.��ȶ�b3� �S��(s8�Q�t.1du�!�|0�}�yh�"V#�r�q�ĩZ�*������M1e*8Y�t>���6cd׮l�	����͈{��Sԋ+si�r��VU�(8�b��
p#��_E֧8j���Y��p�u�V=���ܓz��C�hg�	�$y��;Q .���M$��FOV�����Fv"���]�En�����C�4�ιo�׺N4�qt�1��a��~�T��EZT�]6o�����)�.{�8�q(GL{�˾q&����+��:���G����%����
&+XlxVHYEB    1aef     950�W��,�I�bYa)�9�+~� �*����G�x�Y��:�]�g� ߴ�����͘���盧�����L�7�xFǥ{�q�vv3D;��]	|t��Tc�l
��d�������<)v�N���bC�|��1E5xs�/�nWu涘<����;i MdKԽ��xQ����9l�u�f�6�4����)��b˚sa��7���,�J?z���^5qveYA�x������w���:���O����� �G�v_@Z^ʗ�iyXΓ.	��>�X��"�sA�k�o?�E�#���y^˧rR��P�6�R$J�R������ ���''CB9x��r��� 	�L��"�Q�x�p,�a;�l��D��ߘk����xǓ�i���-�!㤟খ�{�#���0���e!��4�1ph-��{�R�y��N�޶��B���m���n��9���Y���/�/g��)�q���U=C wi�ָ�i��'��T"K>�%X8T�[��Fz��6��%���@�<k�DeO)H܅�4$(�H��ź��e8͞�t��B2���a�ŧ���K��D�v��2|:+X����l������by�_d�����W��I��'R���5XM1eeo��fg��A���ja�ޞ�@Ȁacd��|�-t����6��xz,�d��¯���3`��9y����<`˅������h� bLÍs�̾.V��+� 'J�M�9��;����s�
��dG�'��z��ee;�5D���`�B�'�'A<�����i��U}���J��g��jJs�Ph���?%`R�c���&�.t�Ļ����Gp�e���4��������j���10���u�3CG��oF�MU�:��H��SP֔D��g$V�>�����ZfƜw�_¶.�~W �x�]b� �������U����������$JU(�2h���������|�`����/�-�%A�_�2��cA������i��֞��H�	y����ʃn] )��wV���}}�s��E�6��c盜t0���:J�wl���#i��<�,�����Izn ����)����5�[�a�r�9p��N��J^m���4p�sA)�yV���&��K=�q`=������Hz�u�9��/���I���ߡ���Za)\�X�����wV �6��4{z�n`��$��;�3V����ݕ���F�o��e��Wߦ��IH�x�"�#[�
۴t��,u�	Y=�
S�N)�Pv2�Y��G/��XR�[��|���8h�:����D�xT�U��f`>��Y��@�KЈ\i�➧q�!е[3�x��S�-'_�6�Bz@Ͱn�n��@���D�6a�M�}�ܟ��Wl<��x��md�E6SAԩ��+;�'��c�U���F��S�ejz�����u�Ql��0"6�x���c��%ڱ�Ǘ��3șdP���}���EӑG �T�A���i�K�S�ʃDHu";���u��g`(y_P^��W�a6��(s
|�Ł�Vx�'��,K�ߘu些_�AB5�/�k�H�6�̞�/��Ls��ϼ�	�����K�[�V�Y�rY�̻���=�*�pǕ��̓��7�~pG�7اr��&J`��>���iD"��,�D����.�״�w&'CL��/��_�?/Oّxy�53��Q��q�O�&狽�0����<��o�Y�yF��R�4꽗��|3}�؊q�mJ�_����	���W/w��������6<��v�]��u�.��e"�B^�v�/�KI-�r�k�>��]�|��ҥ�����Ċt`���tB�_g<A��:J�\�,�L��ϡN����ʞ]%+@��f��9z�6?vqK
#�k>����7R(�QLk�{[�ps�����	��V+o��
>=,�T���D�y�G���Zs����TW�vT���~��o3n�W��R��/�fE��H 0,��Wh��y��di�=D�=������`�h�4��>]}�ı$��}6���>#D]&c��G��
���v>yqo�ܻ�o>Q܌P*�8_r���c���
����J���>�tE�MW̨f�R�x�E�Y@P�w�Y"���V��4_\N�Y���^�p��#DYuL�[���Ȫ(��,�a6E����hҔ�uh�mČ6�sv�� F�ՋM�"UN�ۈL�oO�:���f�I+M=���a\��6Ϣ���K���dUU,�-ڰ�>�}�K(Ҩ���b���/�J�B{���5��_p�R�l*s`����\�O�����ۘ�	�[��&:��]-O������� ��rK�>X���