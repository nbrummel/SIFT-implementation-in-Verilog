XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����1��R%%eK.YAp�]�[g9�]N�O'��eM���{��{hf�*q͎�����9t����	Rɛ�V��88S�����>������>ݭ�5�1�.�K�ZnX����U�}�����E�_ý�/�3gIT��FDm0�
#�i���ɕ�_�Pa��?b�O/6�.��/t�P������wbO��?؀��+t�"mk�RG9�A� ���1.�a��YC��`u�gSK;szD�}fa����h���ف-��L}�͊��6Y�7T�+��������=�<�7���3�����rY����a<-<����_{���ψ��--�;eO�(�����{������%qy�ߜ��=�)N�����"L^^�����h�O�0.�Z��4$�K�~�j�9$���lH�Ϋ�\I�be&s�ʏx��ԉ�����Μ���S��]g7�Zj��d�=Ef(�Z���D�;W+uS�o�,�����j{6&�8���O5��,�p�`��6�v�����P��c�����*�,���uB���;�nL��UD$I��ANv?��ojb�TN"/�_Rs`#S���M�su]����<o�ANy��y�\2�u��^��<�?{Q�n�w	�<�LU�GB���=�6e��gn��&j��Ta��·�V��-���:��^���b�s;'hS�5�6] *����v�v~��y���GX-�sG��3&�������V�J��@�52���p����V�p<X^i@��XlxVHYEB    fa00    1790�x	���+��	�5ApiuT�[�Y[P��G�"���%��e��ʪ������u14�W�>��m��B��@����6��S�Z(a~,�9��*��KT�r�M��?`m��ew��B�69"w?���ZV^��hp�f�"B�ip��D��2}2�J�)���=V&�٩�5xT�n�w	(��J摖\l�	"Y���ù	�Q��"���|X<c��o���C���=]�jgD�횢��Pv�,�?�1"+���
&Chl�n�E�>�x������:-GƬ�n�o4��(�Y�]GAH!>_�K�=������@�s?�0�B�̭��t3y�M�%\����@I�I��Y1R(II���ĔA�B��c�ن!!�M��v��b%k^sB��2��#\}$k�=��ѵ��U�'�F�y�B|����7�����-�ς��T��������9c=W0.)TV������j�&����0���a���z���0������{Q��3���Gb�/���t�i(w�OG=`?�bɥă���@<{�E���'��$C�C������%���娌��WT1m0�+��"6�&�U%�xLyL�|�����D+c�tգ}n�S!qP�z@4Db��luꕃ*��;�����;J�l4�5c�hK �-�lY �X�?��x�y�'�c:)̷.)iW�L*�L �ª��3Æ�ׄ���")V�Zp����\NV�MPy�J)`н��PRX,l
hC6W�6w���-�H�׈�N���h�V$ߪG�HA�酿�����/�o1��+Z6����0l��a��7�(���~0�چ-)k������xv�7.�!h��tP�M�f���xL�+�����8@���S��M�ӿa������޶F�Н��L��UaI!��/C͐`14��-��}�V)��{��F�~�d�PX��~��A�x�=��i�Hnjm��f�#J����@���t��M���y`Y��@K�&W(Q��DO�Z?3�[��Pkk�����Y���������U�\׶pf�����I�KHY�VX�9�l��s��m�9���Mͥ����O��� �Pћ,�"������>���� ����9e�`�	��2�d� ֞��)��R(�~ ��o�JBdQ����\8�n��E���N��B���8wP_�����绥(q�̔6Q�� �����3H���[�N)�	Y���uA�M!0��ڈ������!��1��7��zc�0V.`c���>��i?V�(#'�����;. �=�$Eɹ��	��2MH$�֢Ֆ{U�����3���ʃ��S)8j�R�)�����U�sL$uGC/�k@��"n�DQ�[&ɒ��oJ>_�Ko��E��9~���&�Uc߯�轅��`�;tA��z���t�Rzfp�(¬�{"�>�]�/7bT-�*P�������-?��"��poZ���3�n���7�<1��>� "Ӫ�+s���k�j�w���_'�ć�%��y�S���Y#��=/ޥ�\DoR��sђ�:�mk�q;�[���YG,�}��D���w#|OҀ�h}�lEH5��b�a*��ٲ�{�y�qX���I���`G$n���u5�al�6���j,g��8&{�i�j4����5T�e+"n��'�A�
�y�_$���>�Z/=ե��F?D������n�3�����\S�,�x�`��/C�ڊkK�Yj���R~p�y.,���=*A�ʧ��B�b|6�q���hS���\�Ԃ	��ݗ�����k���*����H�,?]�ߪ��z�����Q�O�O)+�����_]IN$51�q�C�1��}�?��@�p�dC�������X3jT�3�;sN�����bK��6��+�-
H� �ռ;~�ɲ\��+�57���xL�>���F�U��.�!����|oC��dR'A�`^6�F��M>�����vs ���Z�����A�1��/\�0[��<���OFy�b��]�*
Z%��<M/�y>��(I1��dش5�R��ڨ{��׊|�F0Nq�a�a�������k�2#3ç�j:����>f1�$��4��?-(���*���ϥ0���\],��砥iY�|^T+�NY�4Cݟ̚m�L��z�Fs`[��$$�48z' v!X����"}�=�ϛ%0������0\ؕ9%����8�¾G��W/�gN�=�=U�a#���`P#�=��;x]�}[� ��܉|yF~l��j	��}
�P�$�68�pǱj{�,�p�h�% ٜW7����F���1�'L�&,�^[S���&
�V�Z;`��F��D>�'	u�l��VF��#�O�l*>ڦ��.+2�V4�ږ�I�,���@˖&��:N�Q�#��*r�t�R�Jqь����a�����xQ�(GK%�u��dk�Ê�ú��0\�Y�M��O�6��F�����|��h^S�s���oݿ
so/O}ϡ�ٓ+�R'XI��
�[QfҊ��YtO��3��O$�#�;�e������"w�@��L��AGУ ���;�)ޚ��i	L�w��>�.�2�jhd��+��h�(F ͏r��o
�������R��aD͟c�I�Q����K@�D�y4op�O�v�G�n!&� ����ɸ��ݘ����X���q@�:)���� ��z�{%�)8oZ���)�p&����������.,YsKI�`���s�T�!L�Խ�\5��bQK�F�����U<���37�7c��S����9�8cPc�?�1����� �)��J:��4��]��m��$h7	�,lւ�Z�K�S����Ũ�i&�f�wM�`Y��sQ���j+��'�!E�çE��'��xY�K��P�!ʢ��tS�)	.8ݠ#(�J!P�Y�u� �x�;}���n��:36E�7?2H*�>z�p�� � ��WJ�^2N��	l�+�:?�T9��\G>q*�&�.��)�ɳ���Z�T�G�o��-�Ø�z��G�D ݘ�{�R���m�*{��[���x\ ���Z���y����go�l`�aU�I"�RP4b��1�$��Rh��i���륈�(X���D���'�����=�(��%}���F���^n�Q8���!�:\�/	�5��g_RBZ��!kꨀr��������'"��/��a����>+���2jZ�����=\Wx�0�r�b��	�������P5]�S��W���gzy�@�� gٰ}��f�G��?��H ]ck��O&�����%`���u[��υ���~�d�q'���t�-������%@êH������vՂخ�.�?0=��E�LV��8�o��G����'�1�~"=�y0{�c�Ow!n��!�0E0E����]�#U�4�L���#�(�k�;���5�D����f�_@C�mJ�Ȋ�K��V7���[�}���X �?:�ɟi,m�0�`1��cz�Ң����}���;�F9 �����������w�nv՛�+�p>���A��C[���<��+��6>I��z幓f��t[I�x9���^�k&���3�w8[yw�8�	��]�_�1���֜ƁVC*�J@��YF�E��D1(=��Q0X�I�ڻ=�v,����h�]��Ɇ�S�,������¥_��ԕLV��dj�2��%����o'#�I^z�(�1����k�MG��nx��d����0x�� �A��q  o�2�뱺�8��jN� h�U2�(e�l���U�$��Nn��>"��\I���{��t㟺`�/WʱS-S�*cg���%�����rZ]�l��L]aa��	m8��=8�7[��nZ������2<�-l�r�ŀ��8�{Ĳ�>�ޠD��ʁIy�Y�YM�� +�/byQ� �gy+<ԶQ��%ǇĀH�j�a�d�Z ��U��S>��چ�;�]��zs��Н"���1x�^�h`�e�{2= ��:������jT0:�(zKY��`�:HfNWQ}���k_Zze;+t8�ĩ҃����!&do|lu��jt|�I �S}�]��D�'T�>�I�H�L�KM �<(k��y4M�lF�J\n;po@�y��N�1���	�7"�R�2��u���<��|���#2����5!c��0T��`ia��gx�ؖ[���@���e��X�#%�e�F�s�ZK��r�Cb���6Y(����p���s�
�@���J���*�ߥ�8����U��8�8FL������Va�ǀ������ڬ�&�N�L�';����`�C�@�J�ʲ/�x߃�G�A����EBb������lp�o*��~#q!#ǁ�z *v�τ��ϕ�z7h���'4=�g�����I���>�s��� Є,�4o�ŔV'
t��+n6��gc�2�:iQr觿�>�T�)��+'��rp�C+Bt��8���2!�\�@&z��C���!w5��T�E��wP� �F�C�/K�ʭB��抨�lz��k�JD��g��ƺ<�SZ.�VR�����l�GF&�����wT��S?IV�@���c���b�=��c8���!���^:G��哃��x���-�p"���t�هѝ ��	��Ǔ�#��C[h>(�,��lI{�ἔe�ݸGa�Gg
U
{�<������2	�q��4U���	&IzͰ�G��U�\��3��ݪ���gq��wݠ��G���U`�
�ͽ�Cͣ:?j2Fmt|�f~�c��lџ�w7z���u��ű�[��I�^|�GiQ(��0X>�8���q��]]�.+�"���\�j ����ti�����}7D����@��|�)�3d6��?X3a-�/��$�>��!4��jމ�7�gň�]zg��ba���Y�cF|�"��"z�Ĕ����.����������F7�E�5��?��M��\?���z%�4��C�	j�?�y���܏���kX�GHaǝ9���#{����^��8-ͤ�M�5�^I'/���H�꼟׭�����Y?�Ft�@^��[�E��F���epq&����y-Bˌ��Q��$��e�X������9�K�"�!\Ay��E@��@P���]�e�mI�N�&��5v��lT3�S߀�r_.��;d�(:�:��ʴ��W�}��2zG_Ձ0
;M�,�^E����R�/�C�K|�(&# �t��tng Ы��|;5d�$J[z~%l���Hmq�N�'����V�YiA:�1:��Zh�4�
�N_��,��	��.����@����*����ц�|ϕ�z#n�ֿ>�V��c�j\WD��ܥ�1:�S}� Ym�VCa��p��/�O�M�N*�CvrX`����8��f�L�B8G��$x�_�ѣ���਀\�]X�������^��:=���JG}ܠT�/y�x`���;�cڎ5xP9w/�W�F|a�����7��cfW��F.�j�jE�^�5z`Q���re7uVG"W&��]���UR(�PR�L'�j��$��c�͢a]%�q�.��b.�3�hv���8n#�5f��������$�4�0��#���+�C�^��g��r>�F+�_�G��ڬ`�qS�"rc@0�2�It+-�,��=�N�|�̳��>l'rf]F��͇�M�}���E��5����1��J�"Н��zGb������w���}���,D������La�N��6�Ԃ�(�M:���X{B`�l�����3�klU�ۦha@�4���z?��|�<�lG��K�y�fv{��3��c�dC�R1M�Ͱ!�:��!�����mbZ07\���P�B7�j4�>��&ʙ5�-7��!6��&h�x.1��q!P��Q����Xchi�}_N��ۨ�tD��wb,�� �g _xA���#���8�9 ;�u�����2�X�CЙ`7�þ=�XlxVHYEB    fa00     5d0���h�<�Wwj�:��V�����3�c�Rz����Z5�/K��V�@?�oW/�`]�6�{a�$қX.����<��f�@Լ�#��/h��k��k� us����F�e�S(\{u���4�� �r�9�Ċ):��'���ᡰ+�p�����}���6��&�� � B�V�7�l9�|��獲Ź��������!�>]�	܂�Kl�xE(�����Mz�"��4n�"�����#-[U���3t�Ģ�R��v��=}�������5��]@���g�R�,Rfv-�����^����hx@e,}�O7YV{��Z�>��,�������vjs������S]R���c�����x7YR��F�#h�X�|��`ɛ��y��hpsmz���c�ι�0�];��+����Ó'�z�I`�
R��`��H| ��Dl��_���'?F�Oh��W�ڔ��D��SIyxt��a��5�l[��'y�*fɏ=ʓW��c��gM]�7�^�����z!��K8❤.@]�C2a�lSw���Cϻ�f�e'k�X\conJj2P����߁�fr��="����x�\#����R	(�mE� �?�.����%!��Q<H�+�s1Y�ɀ�K�f�r����(t�H�?�ԝ�}������lE�YCѤ���-X�K�7�����|#�ǠSu�]yv��*yd�e=��ov�h��O��w�ٓ��&/�����Voc����\�H,j>�G�w�j���ռ� a���-؝o<�A�������EI"P�2E9O-����Z��g���T$J76���7��e��I>EZ�D ]��-J������Rh��{R��������5hN}�D���y��=���`�.ȑ����*\��7g���bS��8��?���O�d�ax�����U,΂������6iԠ;<M�{9��7(��\n��r���^�	I쇥���=�`�_@칝�_TT� ƨ&����P�o�^X��ČG�`���u�S�r�zˍDc's-?���F�)����6�{���f�H�k-��pj�s$���������9�Gj�P��>��Q҆V�aU�k� �7�dp녖O-��`�c���V�f�����^Ar����m�[���ƣ9�'OMu@��� ��")�bu�>��B&C�/�Jhgh(XEi��=�m���D����v��c� �D��)^�#C<ۿ�ȕ�K����0px�&�i��-FH����i��U$�C��A������c��rN�zkG�"��4�}Q�/6�V��=b�i�)�ﵭ��#���3�\����pJ����;~Z���km�ث�v��$/e��ʁ�b�%�<�FM�K>?�+߈�>��Ѻ�M�B,����-[A����u.���bV�/򈦒�d�[�Ih��2�WZ2}����F8}O�(^��#C�TJmeO��~�=��ڣXlxVHYEB    fa00     640*��"�g��$��뤗Ŭ�>/�./��_���g M����]|{�"���sN=C�eN�����ω���mD9&�77B�kV��%����Ua��7���4+>��A���������*.����K�2[�͸�|T���"��P����Se������ �_�0Xʣn���U���p	>ڌ-i-encD�r����+���H��*ļ�9�����fe��{/����#6��%��E*��<r�o9��.����i�uPEn���[Ϳ̄�*� ��@�W�v{b@��Q�ק��|��'㷱�M�Ky�b	��H^ߖu���v�;J��m�I �f��F���6���Pů�]�D&lAh��C6��n�!C�X�d�|������~Úm�$�	c5p:�o�鉧�H�-G�HA0��އ�b`���uDB���j ��V����q�e3�mA�Q#�:'�(yվ���Sl	_�"V��&�S���UP��.a�7��C�3��@�d�VԄ��٠e��0��΂�Ǯ�F�я�ڞ)lܒ2��:�L�,���~z�bE�����Q���U����ΖU�[t��l�U�A�d����O�7VE�T�έ���_o�H��n3�S�*ĥg�!�j���*��d���#����zǯ�P�OS2����X92$��Y�}��T���t������wԪ6N��p�u�'�3\ias��b����
>���O��&�x�
�.������h=2b�äF_�c>n-U� ƣ�v�m	��%	^���O[x���+��F�h�������]��S_�j$]Is����ke���u0��QF�R�k$���>���ܿ�D�	���~Ͼ
U�З��4";~r�j�ܚ����7������������Q�1 ~`y
㼋�D���]�.��%�g�_���ѽ���DD���-�g�v9�����f�V��a>j]PFi����ʿ-=s�9L�;9���>c��JR,K�Y`*e���W:2^QSi>�����!	�d����'C�"��!�T "�[=���b?�el_�y��>��㔼WǏ�F����qϿ��L����;�-Y��>C�f�/5o�F�Z��������
1�d��pq�I$>�~�%�~�A#1�ംF��C��u��W0�p������4�Z�:�ֶ@�e��7�^�;�u$ �Ya���8�r���� ���K:����M 󕔑���_.o���;j_GgZ&�ò�R������V?���?���k��P+��b��Dk��v�c����A�Ge�m�ջ��H���Y2<�*��:���.���������KX��� �0R�[
����[���~\6�F�4���VU����,^r���PEbR��mj;ʦ�gMݘ��i1�&��N��������K�%uG-F��2`��[W�o��ט'��
�� ���i}a`��/D��x�D�������[+H��`�_�B�S�'X�þx(jf�h+wg`ע:������@�����/��;z�Z���F��~����3f(��2���z,@�XlxVHYEB    fa00     5c0B49~�_����<9�BN �4�61��Q���(%F�"��0{�� \�m.�$q�Dc�.J�9�Jf�[8�?�H�[g�X�M;\�n/xm�[=�s|%B���=4L�J�z�	�LE6h���5�I�2���?�:Y�[޾��~^�|�]�hg�k�->��Wuz���>����LB��.q�X���ihN��&�1��Lѡ]�z+HD�{�s��[����e�7��}q
���Ht��SwL~����Ğ�k�N���5����ل��J�6W�F�r�3zV�*���ͅ�\�_	�`
�S��n-o��fw�ux���]m��4ͬf3]��5�*������ @��H���b�9El��������şFXj��Z,`�_�Ϻ}H��4*�v�2�o��13���	΂ad����w2�6y�U���_`��l��lұT�<A�g.���u��>f���� +���#�:3�|�@e)�UJ�'��E�{2J@Y��v��Ic��t���߭8MW��� �I��Z�.k �~�&,��@w4F'FD�C�i�;G_.F�/�4ň�IQ9AL�=�ʑyN�Ŀ?9C0��\}��0^��p?'�Q�����P�[�mv��QZ�Î�U`v�@�
�Z���>|����6�����UO٬ἥ�����֨�� Ζ���3n1M��n�&�������D�|���'���w�8�$w#�6
.?y�,M�@"�$����q����a-`Ɇr��3��wz�T~���e�`\P|�6��ԁ���VM�QbOE��n2i�$�{�4�Z,-��_ʅ8��ߛ��:���+���pi))! !�n9$�-�Ă3���<n!I3D������tM�QG����dp͆Ҧ"���~��=��}@��씍`�ޢF��sa1��lC��s�Ht�I�wU"�[q�G�������t�<�Yó��C�E��zb �&EA�Qץ��KK���E�R��{/� �d�����7��7)��S1*�&U�b� �*�Y�{V9|;��l�4�aS\�S����?1�`m����*�udh�{��%[[w�Ο~C��t���%l�T��]6T�gW�ܙz(�Dy�l��h@�L�'�R�)���8w�����ޱ&�e����l2�zz� 6�z���9����k�?��0��.��Bۇ:�~�eB^���G���n�+���w�p��SC"�B(e/[Pi����<7f�RS9�KP7�� C��8A����5�d5�2�Ϲ�!�[�Mqx��
��J���"����Vi#p�?h?hF���_)�����u[��i�	v��A@mPBgC�IGo�ӹ_7��9:�5Ųn�8���\�;�p�ن�j���x�D�X�kG���o��uI\�@���p�c�h�O����s/塼PQ��h�t�9`Q'�F�T4:�2ֵ�8��m]3'<��5J�XlxVHYEB    d347     a90��~Ҹ��Z%|ƽ�|Af�٢�l�u�opu�eI0g�\A=��gx�GpG$�=$�,% ��}�����j���-�+@���Cs���!��8�z#�V�;:�!i���b��h��p^:��a�� �ӌ*si���G��ދ�A�7V� ��7"M��z�wDD<ǃ�*�!�І���*lJ�:b 6N��O� c�JV��VT�U�
5�/��H~�r,�w�F��B5��B��L_�u<���y��L'�^�h���me@�zmꜭ���-57��u�	�G٩����p@c���x."*Oj��ق�T_����)�����{4n`z�2����0;��%�\�(�Q�Ҝ�kD,����0v�;�h|:���yC�npƷ�8�2�H35"�çA�%&�u�kSDO�;���k!g�Ȥ��ze�%����mJ5��R� P<����
�i��%`�E�1�7uݞ0�M�~	d$�+2�zF[�U���:^�w:�kMEa���*���u�hK>#!.�hV	41� O�*_���"J��!Q��s��5)���
�h,�E����#iaT�݄�:�4��c?�)zsZv-�DCg�Oc[��3d?��(I��>��;7}XIx�s���c8�+�!�/���������}����:C4?�~�;� �= ���tfr⨺�����I�BD⡾��)��P�g�/�D�u��jj�'����v��[O�F�}P��uY,ʬܴv������c/��`S�-���a?Q���������<3��qU	E9`᫗���+�7��Z���Pz"B�/_fY�w�����\���3���<$����Zs�#�KO��&�����&*�&��Rr�jp����������]��V���R��wB�{_>��Q!v��d.<� U����{`����1�[{4*�ǖ�ݐ�� 7�����I���1/}�[Ҧ v| ��ml��Uf{@U�x��n��V��ք�Ww�z���\F
��_2x����Ղ;�3�g�,��DtR�����Ԙ�Ǆd�.i0*�v-2N�w�r�espf,���?��c�zB�>�8�L�bߘd($�Hd/&ڑ�Q�7�D����C�B	�%B�1�N�T�je�oAY�[(�Tj.4�v��\/����g�T�e�ש��*X��A�;$���Mp� �5O�|�s�M�^�_�<_�Q#�qqrqHU�A�_C���=�_�j�i���}ppu_%�/\1g����5�&�@���x���f�\�Ԭ-�<�*\|�#}�^l���p��4�M��d@4����i�( �G�5���j��n\Up�{6�o�wo�;��
���˘����ᶉD2)�j�.��k��w@�ܲ����/7�J���NL6i������VB�Q���^ρ>��U�sQ�$.����,�`dߏ�fwBM$��K*�Oz������]�F<�ø��(��SY�z;��K8��u�)���S��d�:��qE�l��^�v���ݙ�@�Th���Zx��㦼j�X�<�o�|���@ԝ7=�>��L��B���瘭��D��g��l�`��N�rg'<c�4��ʃNU�����O���\߲ F�����⍳�L��S��֬t鋘��oOÒs*#�\r�7�A]��c�J��4��]��>�{_��̾G�~�����Z��cgbШ>7Z&$Z�ttyS�		.��Z�h����	��B`�(�6"��p�Q!EA]���ñ���t��!��"���	�mW�X4t[�S��M�U&äp,�^Ԗ�7R_��Z�ɴ6!�K�3�U�� ���QilJGsz��~"3]ǅ���5���/�8�����b����-���LƝLrl6}�r��z�*�$�e(�ڏߓ�³��g�E�E��?P���������k;!E�`�C��!X�Pr��mū3(�vɉ_�5��{�^�W��~\�%<�8 ��Y7�
2yv?�D���z0�+ 4X^��X�(+���*?�C��vD�]�}Wc	�u$�	�h%s�|%h������%:{�79��(R���ɮ��X>�x����ֈVK��%�\e�Mri+��x-��F��N��WC�`��vv����l7���`��4��k�h�
f�.��%��Լ�a�H�z��	s�*;�F��CC�R^ϣ���W������k~�R�R,�Xk�Jc	���zt@I�%%:;RvF��Ox�� �]~�Ǻ�z?��08��h$��d�/�s��o�1����`nU��o��	���玍2\���9ѨpV�N�� w�L�9=�5��K f��ܲ=?�E��SK�b]�5����L��6d59g?˻�dX�J4yB�NEص;�5���
.��ܶi���"v�)s��Ysf�k��[]����ZY��'H:~�+��5By���RP�L���'â 6�������k��@����b�G���ՠap��M�mڿ�***:zՔ�լ���e��B��%��$5<��M��|�A ����*�*�Ô���B:J�Un3 N	���l�JŢ,AX=!![��A�򁧁�%=hQ���ƒ���Jߕ�ަ�TQkT������y�i�<���l-��T��1~r�c�%�KӔQu\�[&ZD���}	:Y�T�(LfO�G ������$2���J��}ZjL��N�>�