XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���p>�x�"��7��)�n���0��J4�;z���K�N�C!ų�!�q��d��8����J��Ҍ6ک
�G��e�K ¾F�/�b��nX��_���k�d��mqϱS}�HFU�'Ӓ"��.�R{�TѮ�g9�uZܶ��?2������	n��,x��DM/�Y�Sg�Wz9	#��Lj��:��)Sٶ���~$HEb5wW ��o�[�Ն�����%J��K-���P����9��@��9��g�]�7�V~�b:=� !���$��J)�
R	o1� ����ʨjE�_#t�� :����_s[9̩�$~�_�
�]�����!������G�h?��:����5Y`���yFo���B�t�F=8���ƀ M�4�#��}QH��af��U�}�Gb�^�u�h��=M�����2]��S�篃�<JCk��������������W <�;yjg��E��66L�nh��Z��Z�Li�J&F�(!c�����^f�P�ʳP�ԕ�^����� �<��iabg��X'5~����gj�3�	
+�yE�:�V���̧���U"҆��T^"r\�6�	���~��S���yQM�T�~��};�l�؎@�a�������y������g�ճ�G����I�I<����ѵ.�$\b]��uQ���>R(.X��Įh�����"���4�D,0�!P���bp�+b����f�iP��ٞtt2��;�I�����'L(��Ӥ��eQ�]S�WR% ����LXlxVHYEB    fa00    1d70��T�T	&7Ǩ�+�wmţ�n��֩����t�>iI�/�)UM���k>��fH���7H�Wk'%�n�{|��{���߳�ɜm�:�Yx��/(-�"�n>���@b�0BO�u;�
���f�8�rh�0�����́�#y!���}��&�L����H	���T�ً�!����7HS<�� e&�Y��)���F������#Vl.���|Q#�D6���٭/�w���$�1�Oi�؃P�,ph���bq|Wy�֬^+�:\�`�P�Wj�?M�1��F��u���+�`|viV$4�W\n���i���)��3r{�x�\��TW�`�i?+fe�����/S-��V+�!K�qe�����L}���t�^�>��v��ؔ�B`��i��U]�r�N����\��qa+��3�*w#ߧ ��D����d�δV�O�D�����/(�&]�z;���R+C��������@��/�Y���ih�5�]D�.8;L$ɹc��}ad���p�L��kD%ry-{��yp���*D7)V��.�������/j�\]�8�ڧ��}$j[3ς)�� ������Q��t���.�T�3*�K�ez�1��G��潾6�9"LU�5�`A�ī�Ud�����m��TP����g<+�o�3�z��;��p>DZ\ݽ�:i�� V=S�w��b��G�hU�z�BBq�>9�&e���
��h3$���?x(��#x
~:�'I����tt�u�tN*����F��A��+x��hϣqQiA*ll��[�L�lߖ��9��(P������|�� ��JՁzO"OW;9-<�
~�Ay��<�z�_�}ۜ�]1����x�`+�#��7�W0s˴Rɑ��ܻ^ٛ>�,�W�[�;���{�hW+��
gO�M�?�N�sy��#R�f����b���ě��i���L��Jg��*ĻN��͒Y�:��^���al��d������`'!d���4���y��[�?��?��s��0σ���#a9jt�.�ɥ�# �P���.џ��l�T���D_����ېV�zm]:������_PU$v44
�N������9�n&�Y�b2�P�ɓ����AB���d!��Ѵ���u픐`kH,��}o�m��7��enr�.�]�f�U�<����U������A�n�2OmD���+:��`�!fr�5L!�'�V�+� p�����O0&g��t��tP>1%i����(�U6D�a�'c)&�x23��ķj�����\�V>�����2���u���4�)�����z(xc�-薕ф�B�$�p�I9̥
�1��>	�Z��z(q%��W����^��y��Yìl��PD��`������X�9M:)��x��J�Nus��@/^��S�ʟ�ٽ�W�3M��|_�f�����mߒ�k�Wn�6
��X�q2;~L �Z�T!��t3H��Q�6�L�T9�z�A���g���D �%�K�ߑ\&g�i����1چsϱ���i�_�O*��%���K�T6�k �L��,:v�-�}r�U㙶,���U�/��־��ޘb��h�()��7��"et��a�����r0�0�ES-�36���h?�,kE���4�=ȴמ����d~�yT=	;�F�^︈���8�s׆,�)ç [=�)�D�& ���~��j|X���<����&�i������xi�~A[�Jy�K�u1���<�_i���[�rp5��[��� �c���j������/��cU��Β\���.od�e���!�@�N�Wu�@>0S�_�����~<Pҧ��|��pW��d#dHb�~�N�U�{�UR�>�D��c�;*�>��۽�ˡ�\%݄���|�s��.A�$1��A9W���d��:��k��v�A����7������.dd�B��@`�Z��T�	6^Q�3�"At��`o�U�t���=�9�&u5���|�lO)��4X�ɵ�f)�ᮃ�-�������(���>�u����k�O�t���~Nځ��g��]��[��2��C2'�c�����Xf���ku��9j�.�(	�ʟ�����#�<I��7�����:�����'�*e;*�с z�/l����m�t��[�֘C�t����m^9��{,\:8P�`���������c��=�i�9�|�/��'
�`c��Gcģ�(�lU�,�|p  �]�տhRr:
���}0���/�@4����x]�]����b�̘Gϳ�!�O�Zy�ly��)S�1Ο�K�ɠ'��:�4]z����>FʅR�wUj�<��JOi;~�����F��|��f�ַ;b]Gc�� Π�9UXB��q�<�)U+�dIQ�s6�ͺ�]�|	��U<>q��8��C�ѓ}�|��j-�,�"-(z�%p���"4��v����}��y�]�(1EJ9ϖE���~�=����u�T��O�D ��D[
�ig>�06�p�%���]WE#-�R8șph�O��_�jS8��=Rɓʫ�cޡԝ(�Ym�c�0��ߔ4��ؾƕU!Av�jʊ�V8�z�}�Uc09�;��i#��-��Ĥ���T�c���
�X
@����A��y�bhʄ_}�ZYX��b;��E���AmTb��wu�����Y��I�±詞��T�i�S4�i�V܈f�a��H8�H�.U�u�d��j��"V����DR'>t�W�q��J
�*�9s�'3�#G.�$"Œ��:,�c�#ǈ�}�u�8����!E����H+;�[�v��ϛ-�z�������A�,�f�4׃�Tlۤ0�1����Z�jɅ�#�Wgc�s{��x@&Do˾��C2�k�!Pq�om��2��e�P�xJ�#�	�5l$�7!���G1h�)?Y�5Y�bVh�Wbc�����x�:֌�,bB�v�8E�{�L9F��<M�.�3�,C�:;%ph,�H4�IUŚ�"�7��m�����砓�B�tv������t|�����f��k�!O��?���O舉P��+�(o�Ҟ��E��J]��0D��b \ŀN��?>ghAU��({'�Օ�!<��98g�_uUS�m9�]q{Ī6�2�e�e�￭��s��M���:� �B3ױ���ˆ>�赳�'���|b� � ��uM��q�}�ؕGz=�r_��7��2���5%c���D�}� *p����|?ڂ`�O��uy�BtW6�bM��.��-Q1m�3Z�	lKv�	��U��+����������*�ͅ��N��B���_�}�ҭ��)�� �]j)c�옚3/�H��UA�c7�`��%��陣��.�1�r �E����֮�{��dí��M�����
B�R�1+m�f��z`-�&L>��BpEa�
d��cU#�rM�����==0�kAa�����X$�`b0nR��2ڨ�!fYf����B�,�y�T�.�yp����q!�#ѵo��i���j�߰�����djK��U�'�}@��i���'�o� S.4]��[4#а1]����{Y�$PB�+̡�X6$�N�sM��UJn.��s�m
5.C�����.�'��ۯI���[�f�^_�Y~	��Et�?w�A��KuS�;k���������O��"���C�����Ǳ]h%�aq�c������>�8������'s+*�ح��C���;ͧ�ݲ��L��7l��B�r�:,ި=����q}=�)��ěRɨ�f��X{ �RvX
H/ ہ�M�}'����.@�sJ�D���
NS����,R��u����q@��8.�)Ǌt��D��8�2�P�g��ڏ(��F�i��݀_��XЇ������ �K�2o���wֈc����v�C����<�ί��f�=� �&R�]�D����Z`��hy�j�7��
gBO	���2I<�C
D��^�����m0����|s;��*x�^C���!	iJ���Ri�V����␒j�!��ǳ��lqXp�bde��ߚ���|.g�A��)���M�l5�!�_~|�rQ�X��8�(��x��b���Pt\Rm�a�4�S��F��H�����T'9�gB�c�<�k�|61"­[�i���/��=�ы9-��hJ,�����q����7�g a�r�{��e;�nG��	� c���.?�=�����(��;���C{9��F��ĝ�U?o����¶��,��@����Z���I2'��ԋ���wR~:���N��0���_�s.��É��+c_�4o�MG,Z"��A`~9R*H�/�)X��>7Z��Q�+Sr�,���#n0�Å�x�e�������F~��|�V�ɍ�p�,���8�8�k+�GA&�5m�PNuV���{��d���H6���v��ޠ�\����?x. �e��*�ké�N��t��d��<�j0}p4� 4}���i*��'H ww:C���஑s��\u�g#(V�cܡp�O`22��W��ql%�������8~ʆ��N��VuuX ��m����hB1�E=�x�Jy�<|����-�ts2}������k��8�����Kr�y�+D�_����1��QD�U�v�#گ�{��� ���@ΈS���^Q�&(Qp!o��{�H�5�����X�����p��vxr ��2�YjGy�6�Mu���r�'�I5�2�v����!��B	�S.o	���ׂR`֌�q'�L�X����_:˻�C\�"����U:=���}�����2M%I���X��8��	l�QZ��w���]tp�����u������n�4�;	�?��S�Z�A��]yox/GG�<津p�Dq�wHxωtHa?A�gɨRj^������]	�hۏ���v�.\�ΐR����R���H;3oJz��e��/����S�گ`�
t��|��H��C��_���k��zؙ���
N�t�K���������@��o1#�)��kԔ�餹C��!
�������Z��[�����u>�4���~�$�SA��*]6�WI��/�%��� 0����^i�c����(��sJN`�`7�b���S�2)�w���W��/Odo�� 3~��I�.�o�ί�t��Ml�ň��0�7�ۃ�҂,4�������E�g/P'GWbX"Z	H;�@+{��MG��V��������M��τ��n��I�w�.���F"+n�j�����w�0�pk�7r��o��ӮS�AM���I}���!�xj�o�$�d���U��T��4vF۽�9�o~�
dj���emr���
���]�jX(��<����{򦪍�l���Tʛhge%0������8�i���z��PY�@�M�Dct����ֆ/�����{j��'����MZI��u����k����E#����E%g�	�/ꊅ�/�,�8�GD@������Tt�X }�"
 �v��P��g���mX�������+����CF�Ȓ����.(��pՊ�d�O��z�߮Xz/\O����MS�%q����7|���K�d1�/��2{�N�_Q�f��@/ե_|4/i^�N��o,�Ɔ6��Ngݘf7��hm��9��6�6f2���cܑ�:��i@W��G�r�@[���fN����E����0����yy��l��h�)�ߡ�Ԓ/�ݐ�ÕX#����ˏ!�5͘���_k~�Ā?B�2�R`A?D������jA��p���%$��vmP'��k�Ou�[�n��Y���?�^��G�K@E��$�{�Z̘��"���;�G_
�!�jc��j_#�)�����M�I��� ���%~�"h {H�qӰ?UC����4�)�[�ך����)b
Js�Rfi��7���M��"s1�<���x�(Wڀ9K"G�"S���e����˛@��ޏ�W�E�qc�@6�m��,���0;�]ndTH�w�����qJ�h������e
��]L	��Y�&88FO���^ZN�DWg�ges�W����f���B��H�5wH �l/'�M'���G+��5H�#�|Pl���J�J	?�5O>GiDxd
9OvFL�
�>�����z���jdO��_B�'b���&v���3��I�'���C�cS02O-���l�D_s[[�Wh�/|A�z~�<%����*n]�8�v�k9d�9%�R���������3�o� s�/ҝ��cKy �筰T�Vhs���aƊ��D��"������6�u����-1���8.�u6ȕ�4���}0c͸�ڟX�x�4;B/�m�T�� ��!$1��L��2�{;���W�ݽ��R�KwJ*ǂ��\�;/J�@Dx.�5� +����^��m��5S����ݯCm�����}�s&�/uH��O!M�u�����LDkl�=�>9J���j��8<|wG��p���A*�v90���va�a�2�5����+vX-#��j}'�CK�+-s��>	c@���^%P��XY��ʸ�@]]�#�>�?C�z��K\Gr�P��*Y�}�e��u�o�h�(���"ؒ<�����׻2���>߂ͅ��8�o�dFyWe��$�@�D�f�-	x�?+������ŕ1� ��V�E���<����4�$�Qۣ������Pp�A@Ć�IP?�՗��^"���u�����]�C�C��cMb9m�L�-1��J���h�OY���CӢQe�쥹&�m( %��Q3N��>A��¤���N�C��Cp<H���nŷ��+u��"���]	��f`�ӂKsy;z�|�w_�~�p-%��ubL5gl�,��
����|���tel�|'+�办�0�Z�2�b�\�h��/8�MDF,��L|�u�}FA|F��b��8��;����������d8���P�.N��V�ً.*����3���4j��?܁��i�(��O\��@�ζ������SÌN2�KX��W�8t?C@���"�0�<nTQ]��=0�tf�����k?�Ў9��S��X`�"P�-�O�Z��z��-cg�rw��Z&������iF�2��o��NY9����Z�Eڙ3I�)6	n���0�k<2����4p>I�n3�ꙟ�R�FQ��a��k�ǎ�P���Vw�`��ULQ�1�s�*x�#g@04�"�QE�f11�B���op8&k\:���-�3� ����]��"��u��g�.�X���@�~��f*�PƤ$��C)�+�[�2�&x�6�b�m��]J!e��?�xQ��X���	�,��[p~�y�.��2[ݾ����!�� �y�.�qQ���vX�����e����G+�EXa����J��٨�-�<��b�%L��3FDu��Z�N��F2��XA��aÛZR�J�ֽ|`XlxVHYEB    236d     6c0Y�$ �U`����K�|Uo{o[�۸p�I�ϸ��Q���x!(�Š�NZ�'��x��b��Sd��2D��8,Z�lZҒ�C路��bI�)I!(J���d�eyJ(9�j��K$�u=�,RZr�}�u�ѭ7Y�{M��ڏ�B̕<�~X��w���{��>���5�������,8?�\"��W���4�W
N���k�P^(q�)#U�����2�F�W[l{�ח�}�+9k�U�?O����P��g	�i�u3g�<v{�;�S��y�N�g��/̾�u�̊=���k�|_zV0�e^�)D�=��A \^���x.WO5O��!D뵭ݶ�s��o<ڎ�$�T�B!�=�v=6Ex?�[�G������� Ms�'�˯qR�O��DZ��Z������b��E/5p��d;���iz|������M��qq��݅�&���,"lh���3O��� �\��ʐ5�
������
��ۊ.3���\�|!1n���36jn]��A���IC���e��s<��vF\	�E빕BՏ>�I e8d�C�aa2����=Y�Q�hc�2��o!ఌK$�"1��&��HcXE��[�m�{��&|���y�<q>nѤ�X���!�����.�p��9�w�ϙ��wY�:��w]of��r+rh��zv�P2����3���M�ʵ=L|�"�/S�B���>g(�X�T_���Q�c ���l5w��!���3FXGk0�d��L(΄ͭ�/�$�E����Om
��:µ�#�ġ����5IQ�zx���g��f��%L��tȑ��+�ƌ|�O��2)\¸��2X)��m��`}}<L^C��t+��N�=N����8��=�$T�}�v |S��`�����
�sDE�L=3�Q]�L�2��m�t���1W��m�i�S]����M��لlޖE��-�6��yF���X�������>�Y"� p t���`J�f+��@�Yd��?��Y&mX��#l�H\_Y*d����=��B�g�I>�.#�V��Źߌ�V���!H�t8���M���L���AN�x�PD�U{z��<-�*��,�R��δ���/�k�����*+fr�ʞ3�����U���l�񸟯�f��N��їc*���\�����������'
��� x�6W:S�����D<�ѩ��Z�(�IQ�#`�ݎY'zi�T^\�Ȁ(��P���ۊMrI�h��Rus�.gr��-���D���"���9�ֺ�	�1�ɭ��/�8�����t������8��{ ��r�L&	���.1oԣ߱�Y"U�G��!^i}Ue�U�r]�^�k\y{Y�3/x2���j�r��b���О�&���ZZ�(�I5�[C|3��f�����b�zQ�E�s� ��^*�o��,մ����	� A����<�+f�*`�H=0�\�Z�� �����zgy�U�����R�{E�@Zp�Mg,4;*���{%��U����QD�<2}��c�}qDo�E�Ѩ����T㝖�nS
���l���Y��zo)��n�S�׵��GD~W��X��D���a����cmy���Ѷ1� ��.H�%-P�Y�9�;��N67��u/L��&{\̱b��4A쌬rD�Q�����?�Q�.��M������4�?����˭I�\����	l�ɀ���jx����(O�W��O��ߴ�D�