XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����(���OY�d��b�����8�@�U�)m�}�7�Kk�=4<�n�7���N�'���h7t�N0�V�\�QFe�+`��Y�Y@Z��q ���'�ɼe��N�,-|�^�ox>RŽ�Ŝ��-�pL�ș��k&f�b	�KzS��y�ٵi��/���V���"럻��r�eQא2�o�.I�Z��E�{Y0!u�d2��u��z �#��2�m����c7��i��� ��g�?'g�|��5�ا���u6c ��N��Ilk�eϊ�ip�&9������o��(���$�1U��}�_�._0��W?5��-��T����T��h Я��b�W	#@�1+%ʥWO����CB��f�{"���)_K!�[��L��L��^%�Wq���_�s5��`,w+O��dd&�Y[2��k���./e�`�Ӟ<R�t8$,�Z��q���1�=�	y�6���ِ�� 3(:�wh�[,�z ������g��[*_�p�y{>h٬�ut����6Z�`UyH*ͅ��sb@��s-��_�U�|B�N�"%�
Vs�����kf��CvТK�\G1�ع� :$S	\�D���V�s �e����WɛE1pu��Ih#E���1����`�4�\�+�0�u��ێV�	o8��x�ʠ�/�@��������l߫�O�	sӈ��#&=|'��h���M1U��O����֞�p��\0��n�����
"�a<Ŧ:~���`)�2/��:�f�[�q�ģcW%0h���EXlxVHYEB    33bd     c90Į�nI�O�;�s�q��Ŷm�{��m����V�����}w/�_�@nK�"�6�<��P�$���hW,״�gA���m)g�%�t_,��-'r��ϱ��M�V0&��&�,�TΈM�#BA�� /'�<�3������M�IC��v�6'�Rr�VNM���ٷ��_,S�ۅ�8����Ey�F	���KlC �y7��&spIL�,����NR��̾����8�,��0�B(oV�".L����F,��h0��|w����D߬0ށs��b
�R�s�'/S������d�[�$J�ףpmlK���`��I��ڄ1mǭ�^���ѡ+ì�:-BqVsl�7��4a��k(�Gɶ�T+�����u�/ȁ	:m8��~Ri[� ��v=��Z��U��g ��P@q�&rQwm5_��a�۷C�l�٫�k�o�U�����"���Ǖ��ܷ�ݭ̧�ł�����[�!�/�" �� ���/F���%�Ł �k{�y��<ΡR��U�u��T:|ǃ�� �QHI�'�l�~*����U���@J���u��a�@�n*�58���q�^��OS�3�fv	a1�-��3ANQ6o����c�9߃-���Q%��!�O�I���G�4���W	�/Vg�v��d���@s�	�eĦ��@�K9�}X��;�D�YߧU�ƀ"��(l�!H0��=�H�C)&��n^�X�z8o�@,�����ˌz"loG�}	h�N�'X٠x��Z�TH/�1�NH����������3;7�ٟ�qM'��1��˦8��suRB�K� �[��BR(D�>�}�����[��!\~���P>;��a~��V(��|ކ �!�*C���LX���R:�{e��h71�8?/Kv��X7M*f�km���%���^Ͻ�+|���뢊�XR|�2yׄJ��E�ޱK��>�i$)2(H(�|N��?B�&�����HX 0��T�?35��4v&��������;d!�2�a�tB� ˷���ߟDm��rw'�+��=�'�Jd��p��_�k0\����i�o�#[D�r ��܅L>���Ͼ#V�B�I��,���i'�/�5���SjDA{�E�2!np�C!��b/T��x�#�B�d��t�ǙIk7�p0�z��`N�ޔ��T����Vc���֪+�Ni�g��j\y���ݨ d����夽I!8�E7ǜ
����fn�SL�v#�n�M��Z�yáVj�M|���G�]'����!3�a�Q"��h���;h5�p�ϻ��Q�"�>��p�[ Q��N����������3U��t���g)4"Qa�:����4�<qo�Y��	���r���f��yP&b�����Q�8Y$,�(�kQ�0�Q��Gކ����� �Q7 [Wn�,��Y��4�Ls<�GTKV2��N�!�[aX	�7� �94���i�BG�?85`G�	iXT���Ԫ���k_ye▢��lҷGv4·f6��=��&:BHz��4��i�ڡk]�v?q0�G֓���N�BM���a"F�����
ՙ�K���4/�=�BG�SK�>��c�n�B��t��������o<]�̪cOuɏ��FPWV�'���9� [���@��/��m���ˈI30��� �Y@h�=�>?%��rO���!եj�y�G�ؕ_��㛭J�9N2؂�;c�T,��t�"4o&
�R]8�G����$�q��I�	$�^`���l@NX�3\���T$U����W�R��1W�'�)�(\�4�L��+r��?5g��[�\��S��Q����#�M��ށr�ױn�A\a�NiP�tZ����+��[$�oy��/r�t�W�u`�X�Q�;�i+(Tx!:�����y�L��Ê]�<�G
��a����7�;W�s/v��@��K ۨ�Z�گ�(Vc4d� ��x���n���i}��ƹ�&�1S[y>�2K֣ �6���X=)Z֘@�p�&M�3$��e�� T��Y�h����l�wWC���"Y������^,|��R�c���'(rE��=�����ʋL�����w�!��!(�2���� tZ�Q��I�ft��X���I� m~W��$�?����NΞ�/�\L�Z�<�6 ��*�-�hr���W/�ެZ��nAKQKR���	I0}=+LU*y��s+6n�j�������x<ʎ��Y�6�����T�OxF��0��v��_��m��u��s$���7EC��=x'��sϪ�3�
��]����@��8��ux)�^k6-zs�n��-X���o�K�"kLx�Mk^e��R�g:�o���S��y����qA�n��<�Z/�5����Ȏ.&���.�E��dՅp}�Ͱ�K��C{�S۽�Kx�=�.,s�������˫����v�cH���w��'d��/�9��I�T�����h�x���r�ݣ����M�RA����Ɩqq�G�TS;�R0��N��K�eb���C[;�xC%SC�sY�Xc���0+�����>A}���f���"���G���Ra�~i�kK���F��k��������R�K��®7�����O�1n�*acI&����� X��؆���ЇMJ�Y&�GNqz��fQ?X�uR�niй�lI�˒��'���9&����g�^,ź��Žln���l�ʪ&8�Ai�+�V�4�7����G8۞�]X�Dv� �P��'�̞6��bm��vL��`��K�`�����m�,[�&2ub[�(B�|s�3��jǧ�ӂ�nڡR}�V �:����D5�TŤh�=�A�od:6�'
�lc�o�sϮ���f=����:��s�t�*n�c��zg�F�%eN�Z���'��3�ͣ)��W/S�Q�sB��,P���2��l���e�@�O5[9�(�� �?)�H�JJ�b3Xo��*��sOC�<��q0YEQ2�B�<_�!o:~�<���"<&k�_�ec�Ot>�Q�C�����Uղ��L�~�nN6.�孝Ħ�fB@��%�E���=v��R�$��	��m��Jϳ{�Z��u��C�������E�l
�"4$:�-Z��A�Fb�aT?�K�)D�)�����Z	�x0D���/��g�ˠZ{�����P�g�~ǥ�,Ǿ/�:zI?�d��=�)�&