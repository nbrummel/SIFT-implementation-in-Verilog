XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T�Q^�DmL���� 3���<M�}�b��+�hO|��l�C���q�kѥ�������?���*�q,�,Py8��'�(bo�p���_{��T�����{{�陌���Bƙ��lY�;}�C��V �M�9ԓִ��mn{I�S����U�QF�UE�V�8�A�呟�p��]K�S�#o���)u���EB�>dr�C�G|vS]ru�N���Q�U�� �N�q}/�}���CǬlaѝ跇�u��خє��IB���׶5���XX���_4�t텒�����#&��d�hD
4&�JL���Da��P=�i�=\���7����#�A#Ҫc��wF_��w��:zz�ڬSP�ǻ�:}BՀ*sIӵz�cI8��㮰�j��Yc��W�Y����*o s�����>ar(�	��9���ɃhG:*-f�}�Q�[
��f����vk^V���iw�2~SW�y
�l��^:#$�O%M�*8��f�EL�4f�u�g��̂W2�_y��bѪ��s�<�4�a4qk�N-�@��څ#Qq�͇]��L�L=�E&@��CH�iݴ�R�W`�RҲ�a��I��������WƦ2C_�V�a�oay��`����?Z)�ń�C���^�g�hR0W7�.Y�����(�Nc�|�c�]M2�	�kKK�'�*�s�3�~�UI���E�#�A�UG�=��H*p͉B+䵊T�8ϻ��b,Ű�������yE�����&�w���QK*XlxVHYEB    5073    1100�f-���t��ɮSeGJ�V�B3�!�n=�f��HU�jy�&����Z��A�(��7�������Xa���7���4����310��5���*~���䳻�&�B�[�nLl��4He��o �x�(�Jx��f�LGݣ�m�*?��i/�|Z��6�Po���z��S���E�WZ��I� ]-�M��w
��^�Y���ak#��/�>��_.���^[T��2�����E;�q�;�����T=�����O�qV��6vtL��w4��~�qa���o)�7G �.|�`�KFl0�;xR4U�^�5�ż��Sh��QTI���5���,�H�f�T]�61]2�waSҤ �[Y�E�Փ�~�˂眐0��}�����Y��^%{��-��
5�$�k}1���O���a��Hi������rK1�+�e��K>��b֝�T㆔Yhb}D��|�4���OZB����w=��p�3��J�rR@�XJI��c��Bf����P�׉�և�h���w��
�y,��
[�	n͍b}@�WEq�rH���k�����O���]t��W�o��E$�U�r^�����)��:'�!|x%�3 DL�~<k�
�AА��	U�Q�_37<�ί�Xw�f���5�v�J���U7$`xTb����=��}UT1�������$�0�"3�6�X���Mk�Z�?*LG���/.0�ݻp��¾�0������^�W�4G��8� n��@ͦ2~W͊��^V_��`.I��Vr�-f�UZ���}Ƣ��k7�
�W�m�岼*d��Z��/}����4bNto�HރY󰤉&[�>�N�L�Ч�z��C����lP�%�"{��n{�����\Ճ�i��oϻl5�St�pQ�'&b>�wRW�ņ�;%���z����ɿʱ���ο:S���{u�bGH �.����2��y�%N#4YM����������7c�@·�~�]4(p�L���?��!Ѥ(�5�+��2���URwh��/�Ld�Xɠm�+��/ކ_Vs���5"�[}膷2�&�%�}:��;ƫ�D0�&�݁v�
�no�i?�w�=i�G���R�y��|>BK�G��_��� @Z���h}j�L�t�i��`T���ր�#��E��y�ܰ��]����NQ��`m�\��c9� ��+��Ɓf�A�-~��N�=�&�#�?����z�a�x�_��ʲ��~�1��ܸ�@�5(ワMn:�q���j�4�>�ᘩȹk_�{�K�#S�:��� [�PPG*~@����t��(�@a�\��w:P�z�(T7�ҲZ��
�1#�8� 0�y�M܉�"cF(�`QPwF#ш"v�?WrV����j�-�����&�1x
�MU�:�BU��A`T$��9E�fcua?A����ݝ����[���X�U�f+аM��86���qT�BMj�l��z��J���e�z��Z� :�|77���M0|m(N{�"&�������xO�F�o����.n�D��ċ��\�NW��&���L�v�L:yQ���� )�N�N'�F�b������חi瞎Qm�'�^>PB����ڻ�[Yþ
t�V2-h��/�\Q�:�.��Tۊ�|_|�]��/v�/G9��,����	Y�Vi���K?��DLzI�����И��(3 �Miy��=Vw�2��k��Vb�P���:ZG��xR�_J>��-� �t
7��\�\��is�o,C4�=��m[xD�׵��K�����_4qM�J���ߝ���̱��z�e����+)d'���-��~!mae5�_J�L�����6뭑�=����O�^�?���|xj&R*.ʵG�6�^�6Y/�����K��ֺӶ��T����19taNl��=ά��rv�D̜Щʗ���X�?Ij����|V�\4���Θ����[�[\0��W�˄�0rM�ވ�.B���=F�vܬ�5�㻹�+A,�Q���Í��Т�5�!���S��2���>\ԥG��T�g�Opӡ�c��T����;od��iHg?��?6[�R��3G�T� �����\��#�V"�F���L�w�j>�g� c��Jj�,��كdzbm�����B>�zYG�~�ӆ�G3��7�;M1ۯ"���q��|l��Pd;^m���I��b��<笠9�q �o
weC�����ϕ�sی��M�G�J�d�SdX�v��^^<_�^O0��ࢶ��/�����8XV�IQKen��p�F80u2r�Dnt���zN֋$[���l ͩ�q�~Z�{Om=X)y���[���3|w�@�����*�N�k跻t3�9#털;ޒ�]h��~�mq�J�?̈́�w�t2�P�@dZ\�&
��w�o~{��QypQ��Q�J~KΆ��>��kx�ہ#&؄�F��{؟V(=U���k�Ş�=�iRv�=
h=�WO�oE���⩀7t�Ȩ��F"��\�Ǿ��C�m��b�!な�Ld�&(YR���_�{a_Gn��qx�����TQ�)�jP�O������aq��䑩��K�� Ϋ`��L�f�g=���Нe<�3�u@���N�z��h
\&���LQ�Ǔ�˖p��7��C��,<��A�MC���Da�����Q��Ǳ�^��-[�R��|}�Q������	�6l$�^�=������.�D��{>/�A��m�7�ЌM�8��Ïz�������>�u\D#7s��� 8����B\�,���{X��L�{��
(E��fR���J�_�Եq�]V��z~�+��*�y�@����7�Rj>�h�s�c���,�k�c'.��ƭ�nj��*�`��T`p>�K�4{�v�|�FO�3�FY�����m�5�TA9��6��J�1�`�(s[�q�ê1[�g)4�&Z2��h�-Ѝ�9���x���`x;c�q��,~*�ԋw����I�J2��FB����)�
&��d,\˿�������������#/��x��|�����<��I�ʢ�<���&"���f4�6X��6;'�N����\9?N�R6ݣ5��g1��MÂUze��D�<͂�E�%�n��o����6��S�,�i�B&�Q&���4����(�$y|�֡�9�����QZ����u����C���)�i���Vz�1o��p9c\�U���va���7��Vi�7���;�5���F7�=��A��3"�a�'���&�ZRu��`�pq�&L.S�2~�\,�xԜ?�ey�CD8�Hh��%wr�UT��<99��d����DW���^X���h�T�}���\K��i�q!���!*AKۢ�ڡS����,ס}\���Y�~��͐�ayR<S׷���C�����p�wUӅy�Jmus�O���� 6�� 4_�E�,�b$��؇�a}ɛ����X�mH�k9�K����w���^�>|��u���{�k� �� �,�Ҟ�����U�J=R������L���,/f���>81��W���o����#VOn�������0�IҨN��ZЄ�p ���>	�ga������^>?�����j��k4~��s z����?����K�rj��:f�Rf��v�1�]e����t<�Z�l~����7*�Z*�5گfA��X�C���]�7w*���V� ��ǻ7��&;��3ߙ���j��qr؟�|;D����:���D/��|���U3c��z��v��H|�)p�6)�X|�9|O�k�g�(ҙ]wэ�>q\	�����CC�8������������!�0T���1=!�R�ץ�X��]�������H�0�ƃ�7l���?P�e��y�� ���k�v��N���)�.C�O��~��0"DO
X�xq�rT%t�&�u�+%��& ؂���]l�-A�Uqc�U�����I����;`?��mو�
�wq Lr3�jD��q'�X�����!����q?��|��)~�aǃ�%������v;�.Ct��-�N��୸���S���,����?�y�_-E����ӁR狞�?H�ջ�L둈�ĕ��K2U�(#� K�( ���\)��ki�;Z�aW��HX��E��l��( �ܺ�3�zR��+�_#r�i��
�
�M'Q���Ϻ��=�`����Up��|�"��=(�C�G ��@(^�ÔF�+�:����f��iJT��Lt6�LGP@����R�`��9�f~�s+-�ԍ��e �X���DN�k�hE�	����%��AB?�����2�E�+�