XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����"M<^��'��E�)����Ad+���6lt���:c��/#Z_�b1o%���~�\<ҭ�'t��&�{�Ѣ��&>qN��)W�7�DP2���4"3f�!�ڄ��+y��u���~����z;Va�l$��!܉�n9xȤ��,f){��]ے�C�R��%����2j1':;���e�!$2�\�;��z���'�I���b+)�6�Y$��'���'��+<����~a�pa�	TB�?�X��?=�<D�AGD��iĮL�c��,�؅1.��h��
��T���1�Ռe8Ա���b^�j��ˍ*��� ��t���A�f��@��Pj��s�r����}O)���e��g����X��nhBt���A�yQ�G1����@�uf����r塖�����.q�R5u�Kq��N|����LS�x�Q�~���������p_��a0�c�7XQ�i�{�D�q�iΛ��)�3Qӓ�}�c(��4�:�x]�3�LNTB����򖫲k�{FBiu3�f|Ȩ7��p%{-�^�3ͳP§���Z\`%��L�kg،��"|T>�H�����dr�L�iH�V���1��^r��I��]b٭
���"_��6uc��^ �ί*�Hn�޽d?O?�:)9���?��s�{� �O7����3�A�3�@��9ܣ���>��[�*DڪN�ZP��3��`7#��~6��>��F�%���Qx�����{C'+v�b�2��6��1e����]��ZJ����WXlxVHYEB    1427     840y��C必�G�]�Ԏ�EBVg��+�j�	*5���lX��0�r�<;� �
�|��w~���a�����Gj�@��W������DE�����Eop'��z�;J|�W�JJ�o)	�����A�BB��Z1�p��ĐE�?�2�aK!�&�q'+��$"�;?T����xq����ej�6}���&�[�*T�[[���Ю��R�G�t�'�6��k�4�NXG�*?�|"5�y���
��y/sH����� w� �ǂ�@q��	jg\s��L�v�+�*
Lh���@�)�
7�O��k@D��f�4#Z�
�iX��(�g���F+��g{������K��Xa(�Y)vL�Ŝ�?�Q�/rx'��XA	7��
�j�!���|�E{uu٦� '��k�F�y�젓����$䑧����hER���c%,86�b#�����'��iq�Ȋ�l�Q�RF��@.��0�g�L����4v��&2AW�y��Pؔ���9�U���~��34��g+RI_`2w��	v��c��t�W��YQ 2V^�J�љf�k;`��o[�ET6�3Lr9�B��(�Q�fiB��"��\�8w��N��L�Ӂ<.N�/�W���]��!��V>I������#�S�=B;c�܉��A0ڍ���S��hn0�O�3qy�@#^,AiG��Ъ�֥Q��l���&l���Y�W�K�k~#ڡ4������'���Y9Ȅ����&6��l.�(�#�pʶx?,�L:��<�zIp8g�ȅ�$�%k���̙��
�8+Ri�f6e;J�q��
�(~��	������:Wv��aw~�k�!�\�7�@:ss$��U��{.�\<@)w���Uie������ggf&�B鷲K��>��q�6ɒ'��K�?�~4��(L(/X� �v�&�jD|���t�+q���.�w��M��K����#O�9��� ��|�`�������}P#|�=��5�XG����4U���R�t�[����"��9�3P-�YU(�T+Ջ��O��(����،�H*�98Z�n;$m����p�-��VV�_c`-���=��Kl���I���IF}=��G9̹��I������am܉� �R,0�Q߁��,��6�Y��a�g2^�>͔qg�pz)���L� F�#����+��S�w,}��%����q�O�6�,�^d��&&�U�D �hA�$�?�KH!�́J����c�`�{�VI;��òţN�sx���!���e���RW���H��3�A����'�ؕ !�I�0�yCR�[�GU�S�}Z�#ЮbP.=~����W'RL��^��p���`V=��b�kDq��t���R�q`���)�ς���Sgz�]f�VS����)�o`Yn�=��cb*�QBD+����!���^^�f�jA��a-���d���3}~���Xi�lI��sN�-�_��xw��TG�զ~�t���V N��Ր���zK�j�<�4��ɽ��Սǂ�#T�p�!�����z�H��aR�9�H��� �G9���������A������`i�z\/��Hc7���l���EB�Z6;)|/�L��+u�(�?^��Y�w�r�t�҃���6�}�Ց�®d��%���*������W�8~{x�@�9Ѝx�2KZ���|l�T�����r���"gT���}8�BP�2����o.9�rG��T2��w���m�����Q��&�����dS��,($�5����a��#ۅJ��h�٧:b��`��\�3�9Ul��b�7����{�-d�F/(��$\��8+4��̯'�\B��1@&c&�v����&����r�\;m���>X��Ĵ�!� �kEvB�a�86�FN��� �u�	���kG��Y�n,:?���w|�*f���:�6fdm��д &�ey8Z1�ױ���N�x���'td)'{��	��6�����~>�b�&n��Q׶�ٌ��q���:�=�%��.p9!��ٸh��@e<�o(Y�)���.x��b4���ߚr�u%����5>��S�ֻ�aOh5�.�	�ka����kk�/q���QM3�������wz