XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���`ƪ���^a�?qB;'^Bx�`b�]^|�|�D��9�>��a�J_�SG�4��*�p칉�Q��e�&x�9�lu�]�sq���"�~��2Ц�2%VM՘�+�fqVB$��*��*[.����N��	�=�b�ʄ=ĊP��6~�gX\}��r�`����$`�n�I�!=��N�]���'p3$��j`��8�,�rI0�y.�U�J�$���� ���Cs��d %b��b��1a߻7��1��]��,6��3n���\�ҀK�ވ�C4u� �K���m���'dpVM�l��?�"�'�wr�LW�0�IxO���ў�pvGL�U+$�΄�,!J�����3o�aT��\״-�ѧ��L?׿cm���^C����`�.�OnF��O碫W�x1��+-ߕ]�lkP���\�����An���Jҡ�A̘�l� Ec�����GT��'Vߐ�O�p۴C�)�ӥld��45Y�0�[����(IM͝��`+�fT���ǏT2��-x���I3b]������Dۖ��i1
���b����jx*����V-��.��7�":�/#���$D�"k��՗����k�����h�P��ص��#vM�x	MF|��8�	K�Psj�%���.}�,4��nz]��CK�I��h��jS,Z��d���|�q�1b���'��ɧD2:�^9X�dg[Y!JbȌ���K:�FQ��K�V��~��t�a�g��S�p��^DXlxVHYEB    c6d9    25d0�g�\� �1c+�O��l�F���"Qo	H�_�1���{BsR/���fK :R.���a	#�5{�����"u��C*��\��T�P��=�F�@\��:�9�V�Ԑ�~���B��#��%(�ɌE��� [�;4u�"��t���X�b��Qǒ�j� s��q�W;eL5�����z4<<A��x[��Q?��;G¾
�0YD��nїGɼj�j�v������h����N.�*	mC��A�$:��7���yrJ;�����ڊ���\.[�{k��-���+/�������@���x33uL�BR���a'*�����l��w��y��Ǖ����h,e�y9��#�
��sA�±i�c�Y	��_�ן:��C<0�#�e���pp�}�b�1K39���6���u&���;GGcd{J�(���5�N*!!� 4�
\b��wBQ��W�c���i������UV��0r_/��:Z��Q����ؑ�/��{��)�b��yL�ُRɽG �ml�z(��F�F��XZN���jN��($?�H�T;}=���{Кo�� X�mYe�i�Dv�>��W�?��6�R,;e�>�A;E�S�t`�qZ¼���˷�����b�N��2/xW�%Ƕ�^~0�^���iJ��cq,dd7#���J����pt]>��l]�_��V����7#^�O��
o��$�дK�2� �[�����n��wV N�B�(;3<[�u�)��``}���+)-P`J�.�ۦZ���N����6`̖��g����nY��Qz-��br�3��#�Z�2�%T੬B`�nÔf��+_�p=�؊֮����еA��6�o!�lG+R��!���nw�*ҁ�4\�dv�d+������xá�.�D�j� �ѩ��k����g�W�����H���egS>���8S�i�LC-��Č���0>#Pg�Ge�X��\(?�X�E����d����˧Q��(7������ T��&IwA��hej^P�6{�w���.ȷ��1��Z��r�A+�]��㝙$L�J7�3��=���zzet��R�� r��D�+O)ڮ"��*�2jP�˲�]~̇���^�K����)Y�i���/��t̰���� ��y/�H�}|�i{�;�7�J(�ȞlKH�����>�ՍM;��*��4P�T~8Թ�J�/'��p��f���]' "^�@Ȧ�#���ʿ	z�  .�{�OU/�N�����L��4���Gle�"p�ԋ�irJ#5�"�b�q����ђE���V+-��hC�����J<�З`�?Z���]nY8��|�����	}P.�����B�@ɩzpt��*̻�@��V�z˻�dn�W��̓O�'W��VJ�T%\<k<T�0X��=��X����N����)wUp����04���ۮx�G�p@����>��[��؂^�D!�Y_��F�K���e�8����f�A{����#���&�	W4������Q�m�����X��N���;3J�c_��L��ҴL�9����S;�S>�\��n���Ræ���4���m��m�a+����4X���P%9/ɻ�%���"�K���I͍����H�AeHC������e��3g)l�f] �v-��(.�8��)���EO;Q�0��XC����XIPZ�3�
舊�e#�ja�X+(-^0�'u��,�Z�O��`ɖ�$�� ٨(y�8�m���n��G��_��<�T�I��e�xD�3X)�I`��Us H�o��b�tKYBsk�b���A��)ֶ��Վ'��Xm�H8�@$gFc-���].<M�I��8L7ɵ�o�|b�!#s��⽷)�D̛��p��Aa�(�)������斖�����'�쎣V'nZ�WP�2�q������G��S�Z����^h��CA�u�n3}���<o�а8A:}�h`Rk�AE2�j���䝿i.�h�E?[�|�e���������Dnk�;���׽�X��������U��c�L�&J0<2NyZ�I.lKI����.�6�g����7����V��/+|60�^k��^5�D|	(ǠWRoӘ�^�L��y;��;�]X4���ӝIB�I���f�e�8�:$)��r"^�ʫ�����d� (��+'��r��V�����&n{*��J#�f��⁾�O�S?������5���K�v�rx���I;`��t���n),�{��m���E9��x��HI���Y�*F�R�{���}D�O���`|����cb٢�7��I�Fq�b9��=]�;$A3	U��;/�ʶѵ�ycQ�W�Y�����W�M�.���W	�pՄd0K����6y>��� z��Ԡ��_
����g7͑Y�ﱶ��`���z���PHIF��������t��?��x�����%�9��j��#�"yV��P�Ŏ�����,����]gșNP��� x���%��h��F��<?|��l�#R 5R��`�%���C��Pl/�0���Zr����8�Hy<=L	�s����!�M7):ǌ���&R����/�T��!{s�M-�1���E��2�z�}�-� �
�_��_&ނd��t�N��@_�	���ʹg�0�<k|4�tX:�(�֗�h���X~���!�ZR�_�W�k�e>6�o}@�p͂Y(Ds�S�T�QwlB�Rg&�@7��V.x�)�)�[�=�ZN�x��!ؤ�����y�r��k��4�M����69ҕ��̆���]=�@}��y�M��K8���I9��ESU�����:V�����)��CR�R~(6����=.��e~.������N�צݠ��Z��#EI����K<����6p8Ns�v�(�4}��u7�`���H�9��#��.T��l���%��2oS ��}g���(x�fbP��f�s�.�T�w:Mw���֛y��\��*"���_I8�u�5/Ba��)1j:t}��h��9�j����~���v/�eyc��U5_�~�;XI�8��"��D����(!\[�>��d���"v+� �7����[�0���r�h<�6T���:�L�Q�<���-�����ߟ5��΢��^��d�b�X5�� ��~6�����F�����*��@8�.�]9���G��k2�;M�ˎ(�!�І)�G�;<h	�W`�Aj͇��>B�d���;� _~�@τ�Ck�Z��T�dz��:����E����t�W�zÍc��s�8�:�6]��ݛ�Ae���x&9p�$�C��aK��	LT����n�ҕ0J��"E&�BX�;�a?u�q��!昮'C ���i�Q�x:�m����l�l�Ӣ�x17lQ�r�	ay��ј=,L2�tT(�$`���Bt�rGȀ[<Y��.����t�)�&����mp1B�I���0��޹�X���-M� Q�U���.yb�{���)�qQL}K�|�����۝"Qh�e��ϺK��%TbqS�;�?��KHi�I��ш:��~CTc2dK�If��W}b4�!R��-��i����h��8v�;C�<�A�!�ڭ�oM�	��#6�\�/��|!Ă��~*2iS˿Z�d2��J<�S��hq�9a)v�Z�*���dޚ�{���Y}�GRg��3}��*��L7�+��6�ٿE7m�9ؕ����=��x�;�*ȍ��n���6�W\���+�"R;ƀ�-s6�����(��s����ã�b�$}�  ��'��B:��C���ȡ}:u�ʦ�)}>��~;��/�B��\0��
ꑏʻB��O�d�c���E�y�K�;�IJd���!#@^z�r^�I�Ƒԙ	ޙҊc�C�0db�JF����Ы�)�gy�(!cmh�2��Ɲ�ha���J�'z6�g��>6�`�$dq�[Q�3���+f9�����]S��C��ofb���Y�����M:X�N����!'�����)�*Q�6�ypxu@�:�A�@ʡ�w��mf�{t�R��ɪ�c���:�dh����9������ �̖ ��.���v�O��t�X��yӑomN��;�ˎ8�	fܿ\|�h1$P;���w���+�6��}�\E�o䗖�b:
	�S@��rP����>V%Q�<��3�(�����;��	z�a٘�z���!�F���_V�9 @0�T�|�!��,DP�)^��`�!��Q����a�� 4��#>��\A(sT���O%Z2p�)Q*B�L �(����A>����o���0�-���]�@	4U�Ҽ�v6-؀3C}��dLQS"��ݑ>�y��	Ź�1X��
a�m%DAt�Ӳc~����:�����^9�9�5�2���j�Ck�8.�y���('ɂ�s�	��I�vla(l��@�e��đ��7M`!�#��XR�V 
�V���G~��6�{�[�B^),{5�3f���������_�1g��~�o{_�iq��CXG��ƥX�����4��Ki-WZԯ�@��֫����Z&�ss^ ��Y�q����m�8�ƶ)ӛ1ͻ`!A�H=�L5��7�E�7�+E� ��$<�䩬D�A�9-5h��D�b��I�������5%}�)BN냱bg������D�}#���af�*+�,���"��(&մ��Ոm�~$"Y�k��+ՖJ��p��O	�8�L,pٕ�PVMb{-���֩S�s\�7B�����ܞه�ԍ��5���z��r�`��њ0�SH�B/�yN�iM^�%W$�����d�m�5��&�o������`?�����|D����͚��"Qv��	�i\��@��ug���l�@Į�~�#�p*"�t� ����ؒj��Y�������M"������&k�M>��\)��x���Hp���z�)�@'�͌ү�2J5>�Gˁ!^g*�������H����w�ȼ���8�o�\(b�A�� ߑ�D����ޛ}���}�B�ª�}����|ׯ�ڏ�y'���-B��l��~�����݅
�s�-F����3r�V�.�?�?�����ԍ@C��H{~Ë�D�2�y���<�R ���P.]:@b>v�4Fs��\�9���;O5@������>s�	����+��6�T�7k�����@��$
�W �mWZ	����<' i�?�Wqie)�|���F�W�!'"���V� >0x��X��ڔ�Ybn�/@����)��V:�X*w���6��h�"װ��:�\�~^�p06;=!2��~ړ<�$I6)Wޔй����T0ͱU��A6�셪�9x �(�O�ʘ��3(��6�".�i�� �hJ-��~���.������ ��Ѳt��U��,���C`j%�Ó�+c�))�NL�5�������,� F/�jg;�9�Տ��g���O����g�Wg6�C�K�	�����H�y����D�u���������k҆��d|ܫL;�>�%�̓�@`VZN�}�2�A60!N�$[-�Cb��X�֤/�Sv~��M腦ٻ)��e
��ϳ*E�l��v�v��C�>���W�%U;J��2���(Se��d l��_A㖛�h.\xw|��O-HD/�i���	<[��~���G����=��DG>og�-�>hA��i�U���(n�z�L��k��Εje|�"�ոV漮*��|do,!�[�CjP9�U�zȏԸ�k�X�(2�i�ȟ��y�т�~�"�<SW]"2�B�Cgݪi^�a��2����%�w��3�z�0-����Ro��l����n%d��~oP��n��c�6�Ƽ�N!�M���J�]�

�����`��#)ZܜD2�c��Y���=~�jE���kA[΄B-w���e-�nq-i?�� ����IW���6�\��NF��ZӀ�Xm��*�%z��1Tz ����6�d-&�h\�"�k�=��P�$p�JWl�-F^l�b��e�ѧ�ȳP���|�N)�M=~�5C�%�[����S�q'�5��Տ�1��Ӿ��T�6�v	k�׳G��Һ��4���<�A��1�C�ayo�ӆޝD���j~\�2�����f�B�[C?ɳK�{�R�??V������2L��,3��
�+I�5�*�	�� ����t'��#N�2�xi�W��&&���=+f�0�a$���*�=�$j/_���!?�����z���0~��5TS>�Ȇ(�@���69��:�{�U)���q�h�Ȅ�ZQ��d\��������%#mBRŎ؝͗U�vпF���z������]F;|����^A�an�~z�#�-�2���_k$Qk&0E�)��H*��������_���2����&�,��$c�`�O���U��\W���/s���4NS?;ʡ���;�@Mo(�y�q�����m�ñcL���`j��|����͘$9��\zn�J�[CKH �8� ŏT-�I� k���ljo 3*�j��B_~;c�C~��ͱ��MPW����)�A����!�����ko�l�\���ԯDC;T�9#��c���5�dmb-gwܧ5}8\��x�U��3���{�w��l�é6x�¥J�"Y�_4XA�vY�+S����w��$�򋄶7����k${SOo�V���X(��9���Lh]K&~ߢ�[[gL�#�v8:�����D�+ɜ)b䩑9�x��)K��%��~Bk�Ն��vqyo9UM����`T��UXʣ�8{�oUĹgDȋӝM� ɳg�=3c*�?��0�����}�ø>�����Ň%�Kj�ƚ��X�KzW�U��}>O|Pz>�ބ��T����d��^	SW����7>;8�y�y�������\FQ���-,��r5w�"���Ἴ$Q���ѲM-����g�d��p�M��ܚM���|ҩ�1���!J�Y�*l��!v�Xp��F�壵�C� 0$C�I^��F��*��B�\���g���c���&|�g^����jkDF�x1�S���:X+&cS�[�Bb�cR�m+V���q��?^��v��!�N�#�D�_#%��j	_�4�bO���Q��rP�ݒ&�[5���U|��5�k���!>��&f�Aq:{��� ?� �&jȻr��.�6�����v�@̫�_>���+,�׋Y��=� � ���
..�����N%�{G+����5�D���9��A3��Q�i�{x�8cR��j6�<F�B��V��D	1	'����7�&���Q����|�j��9�{�GķǄg���M��(�_y �*0� WB
�%�S���0L��+ݼ����9���j��s����pĽ'x��Y���N2;E��]J�%�����U����#��Џ�uSDa\�0&ߣ��hſ� �:�f�e��`:�b�\q� �P��}k��]L��XsW��g7�Z�W14�7��y�B6���[���km�Z�iҊ�0�lIv��߂����ƭ[�[o�Z(is)��x�.�5��Eb"���uΩ/�U�|�����SY��}�������шF켘^p��9�kD�/�h��K���牥G
�g��}[����Ra{�����?��✲���A��=n3��Ym f.+���e�������B(}_K�B"�x�[���H����vP j��[���Y���~i�ґ��%��*,� ��֧�^b#�	�(�KU����+#CͿ�J��u��w��ʸ���*����JeՏ��E�-�i]%�ŐW1=�g<������:��su k���ŵ���C�
�Ӝ\��0<�lzܙ
��
��x�-rڅ�q�P�~��;���?��㻒���V=ӿ������O�\�[�������;V���-w��ZE=�X�E:1x����zj�]�5�}/i�Cf�� "f�£9�0	�O��ԯ�m3�w]d�'�l�����x��U����o�纫�P�^i?n)���?iۨ����<)MVH�}]��^�0S�%��>Y�۟哰��� -����{��|�$C�'���"S#�X/5��s�&^����d��q�\�y�?M�����[J��`|�ȋ���A��=p���"���3�q�pȓ%畊U�/Gc�֣T{!���!�=u?��֯8k��u% ;/�l�
���7�es�ϫ�_}6m�C㧲l@Ɛy�8?bR��Ƿ��!i:��=3�	$����c�fYI����u��\BY���vC��o� �����m�+�;[T�-$���nOr��Æ�H*\vR�8�c j0�`�9#��ȑ�R2��jUn�2?岘;^y�	��z�۾��s�[֜�89|p�{�Nx���p�q"�[���$M��d��N���� �Ly-��.J�X����
�J�u.Hku���Q�]޺BG�MtMώo�vS\5KC����w"�u>�Q:�y��O�uz-žZ���
��KXy�@`�ݛġ�4R1]�b��a����q������<��.�5D0m#�U��'��"�fIh���7~^׳aD��ct���Ljј���[Y�����������1�~��B��9~�ʀs���łlv�]F4�z_�5�6�v�36w�v�O��\(��S��.��f�$*3��X��舆�VE- 6�L�B<׀����BJ䟊ŐK�WN�~cuv�ڊ�V�#���ӝ���Þ+ �/@�f��l�\���7���l��n�a�w7�����̠�&j5�f�:l;�e�^���a�_��:���8��*8��U�Y�c��zw~�/W� 5�ep���Ǥ+H}�b�-�?��F���|S�T��
Z��ts�QBP����o>�nS?f]��+@�U�V;R�]��t����9=PL�X��)�/�6/p�{�Un:^��д2���u�^ؿ��˪5���\��N�d��2�D�g:��m�r�3:�c;qHʕ)��>�
��W�L�:g�����í��X��j%{�3wKP�=��G?C��Χ�[	7�7�[�Wx*�nr�-*�~�㷌��hģ��ڋO��gN��ˌ���h��3�T����h�øm*���+���WS1�N�p��]�&e`fvb��]s�Z��$��Z��r����5eT���>+s��҂,�Xi�c���?�m(�P�j��J�ĩ<����K��6>F��?Σ��U^��(�.|{'��޺�a�-������h��Q<��Z◯>���}�9��>෋�a�&bts����"9�޺��A½v�^����U%������k�߀>(T�����U$A	{��}>b�Q�D��+n�9�7b�)6��3�w�׺lVoD?�8�� �@�i3��=�UJ%�w�AZm��}��%�5��l��F���
�莙��'�A������� �����<v���>��r3jI���@d"\�0�#�����*�X-�/+��Z�Æ1��{��
���k���h$������iכP1��`5n��lŌ�j?UD��MW!حX��!���L�� ;�-���],�)�׈���:�dE�J�