XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��f&�^�H�Yr�=��cِ*h�I˸
�};�!�\��s��	�����]�GCfcvW��"���B#j�@m��(nMf�v�����k�C�Cs7�<fِ�;��RX$X�&�x���|XD����{��Z%���%�NÿF>�J������m@�n��޲>C�_��M��i��w��'��������4|_�u.�񢗿��@��rM6d���%e���H\�C-�ݹ0Yw�
�º9p<(�#^NG�_Dz��{�g&�.b	��2���9���.�x~�f�C����_����3�P���ޥ��,�q�����������z� ��?��>t��DO�^>��	O_�뤴�ne�A�I椨
A���4�)��6��+��E�0c��LD�'eL��ُ\�ÕP�� �O��3(�9d�8��]��'�]*J�q�Z��񥌑�F�a�@����r�W|/�yl��'	��5H�Co.ݮ*�|���M�!��|�[��P�9R9�p�gx�~F�6�qmD	@��'CQfT�t����,J�."�/[�T�F��`K�{��݀w{s�#��n`/W�v	"�A�I�����8���.
B����"��O����k+V�W5A�,�{Q��io��L�X��)�p�	�I$&���T̼��P�o�ޕѲ{D�w)��&��|�mx�K��S=P���6�S��[� O��0�fjl�����)���w��/��g������LP�|i�lZx��=�XlxVHYEB    fa00    1f70MO�Ѿ ��]0�bI��W���l���1��\�%���y6#��Úw��i$���]v���!]���j�?����ȑ�=����6C�b��A��K�i�#&"ɏ\#+��������'rd�	@�%��$��_�IVi>����Ͼ���P��n��ʪ�>߭�\� 0y�y�8�O�!�|3(��āVp�B�俥���FHq\^5�L�S��쫇��V��xB��;�G���4�1���e����^���ks�����+($�*�c������U�����}�����Ν�m���!q�/��uV�FĶƊ�Ta#J�W~9$��gA�"���Hc������F�[~�f��k5��-������d�_��l�	NW�0������	Բ8�d��o+�D�8�iE ��u�x����+4�^Џ�80c��*�o^[;G�X�a����F������~r&9�ox�Ш����>IF�*�J�S���x��q�� �(A[���Ǣ��"����U_�nf$��*�&��ur�^_���w�t�1~�����hC9���v��)s Z�� =#ٳ����
q �f˹�/u@�X�  "y
�I�����jq��
�jI ��	#�?���Z�	���X����[��WեOЬ��-�"�7g�C�厊%���x�cQoh����/ߎ�������Nj�E����"�>*�T��MTi���tYC�ǁ]����H?���>h��LPoӛ�6���Klh���u�%]�E����Ʈ�{`���ؒ�)�;td�<�_��ϻ��99��p���(eN y5�|�e��u�v/��f��4̜�����Dwc#M�	�dE��!Z���*A����0V\�w�~o�ȩ����2v6��i4�X������b9�"A��f�֞/�\�Tuw�	7l<S���5�y�Lئ�O�
1�Z�Y���l`�o5��E�[�1�-*����x�l0�?�nCp��^	�EE�&ѕ~��/�c�=�^]����U�(w�k·>��8�SE�5rUV��y<�©i�$��p�u�)H,t���л�8�=Bjxv��<֩%���^�JF<�L{:��ɽ�1>kw�\t�������g�@	Ɇ�B��|!��ӄ�V�!a��k��Wd<��pt�	M�Ҿ�n�����b� ���V�C�Ef|�����q�?��<��Uy�Q~~ů��U�/��3��l��>�����uѽU.��F�?u n�2F�j��=�t|:[�LOWJ��f�Ԗ�)z����ͩ�^�l�v��I rh�5!�*Le�qS��Ɏ^fB�b��'��u�!���h�����j(��#[����_6�F'�|	TϪ��_]F V[$���_�H:���5�ZIB�E@�wIs&Y���������F�ʼ[ׇz�5?<�Qͺ�b:G�n|\O�_`w���ﾷ(\�r:���rh�qV]����-x$7D����f7k��}��c�aԔ�^fm2��L�����\χ��5�afW�Љ^+�F�F� �$�VF��.é���y�6l�Ϡm?.�6�������i��ʢ��T�C#'6f��k��{c�>ⶥ�a���|�-ʋ��r:�0�/M���O�qb���=nN��cV�	d�����_^:h��uP����R ���ΰ,X�4����sFY{���T�w͒oit�!)H�����vѥl{�k�x$^�GP�j��-��Atݍ�F��H�wΡ�]�MD��G�k��H>5�f�����IO7g���X�t�=��Δ&E����.�i�ppb܅$8d��m�u��ֺ������/Q��M�������(&j(c�<\Q� �(wC���Rsv3�c��V���x��4�ݪ�*�U�������㛲4��;D�������Fx oP9�PP�Ӻ���$�z��\k��)R�v@g&��ĝD�@v��n�HY�`��C��3�q�[���8��oY�Q;?�!�D}�E5�]�ڳ�X���h���I#� '�G�N��ک������\ 瞞��ҸU�G
��[��T�������������eE)p�[�@��)����g7�?��[|Ҽ~�u���!w�c{��}�!�c��[Z�d�u�=� �i}��I�ߌs���#�Z�I��aj���TL�]o�"-��z�k����uE�0t����'�����?��(9��=��XO?��E�h0���d�P�Ps��S��$�	��]{$��TU�8���@�v�9Bs���O�sJl�x,<9�����Jx�d��b�>r�<���m��o�BN[{rcQ�]�* �9r�.=7gu^Gl��}凁��.kQ�Є��F#�!��D%���"�T�X��1�! ����i.fU�\�L�=�����yo0�e�l3$�RwP�G "���lkX���p��F�pzc���������E��(Ex���芸�������.8�z���յ��CP���QK�l��U�s]478��f����Mt�N���!� 
[����G��1���Iҳ7B,��O/�a<���B��~������ڗ�k��3����m�����X�&����'�X�x�?Y����̉�`�2*����w>�����)��+�G�3L%n\�	q�8��h9��~�f(�NaW�6�iM#�>�4�����z��$ψS�3F��o�.a��93�N��]�0^�m�(E�Œ?����}��0 ��&mp땳�ʺ�|(�a4Z�1{���%�����s��q�+D��E��Ǡ)D�k�>9aM���;�9�_ ���ϧV�&N����@�r�ht��UbL`��@\{�N[s�B�@�E��E�-����$a�	�A�=���]RI�.����1�wO�k���z֡o?�B��|���JQ`�����U���8��G������[���-A���|��.U��`~��3cɱ.�+D�#s��[;ҫVN��s̿��Q�I&���l�@�zl��(�������U���rS`���Ջ<�d���R܄���Ce2�([&�W��l�%�U4�����Z��
�;�d�dr�.mޮچ�ŮV;)-���������#�ȏcP��1Q�!�%�/�� ���� d�1A�Y��џ�b��2ro��+�۱AXd�h8=������~�T��M����MKxr@{�-l�}�?з�q=��m���&5*�6Y�u{G���$�:�Lѥ�l<s���"O��͖�1�������ސ{?!���쪡��e_.4��^����	�����T-#����
[�
isE����-����� >0O�^uw��{J��Ĳ/�z�\*I:�{�L���@k/@ܑ%oc*�Q!����}�d��PȞ���*�ي�w-����v��W<ޜ�ȸ��P}���JH#Ͱ ��H�1��E�������R��~�4���|��Z��ɤ�bН�z[��p�����J��K#���q��ĞՂN>Uf��\>t��5����Q�W�Ծ�pN�:jO�/��mS�f��y�1��m]}���T�M�:č��0���TC���E�EI��IݭM�X�uV���@�n��3�Jn���J����Y�U�=ʼ�����m �S\	���D�B�n�B����R�G/�˻�/�v��N�P����S$�$�@�G>�]��v�����=q�f"�����;֋�|�V��j9
�aQW�M�k zG!q=�O�N�fӪwò����
��v񌟽��.��N\ï�5�gʤ�s��01�G��=M�x%=�(�|xt_ �\f�$?�w3��w>�
L��,�����0���Of�����Vg����{� ��/��
䎖�Z�p�m�
�b�}7���)D�� ��n����]�:��Q�챍��7X�G�q�i�2��G���x�۽x�~p�㺞=�vp��:�ԃ|�����{K��`���{�̠g�wa���40\�"� _b̉)��E&]��[?м9JF�0+*��|q�|?��C0�<�O���(�nl��#]�}T��ZO�s�ᠨ��ƃ�������v;�]Y�"Ϡ�<$ڭ�?dT��(`&U�2{�?s������;+�T�Q$ +��5�+��5��O� �M֢a�YI��B��	�+���~?_�_�(ĕ�ɒX���Ej��/��S[i�U&(�О���)����pT�e.F֠]I�rxA��ƴ�}�	���'<����t����ZE�b��WQ4sV�Q$y?��2�Գt(y�U�_s����LI���MM��H!^�6$�k[�7:(�-��4��]fO������9!�g�)�@��҆��` �?�2��k�c�\$���A���y��7{/u��.�7����r3`��v1VN��`��RmD��wxڻ������5!;����uL�TK
�� ��C
��E�To�G��F���N��n6ʠ��H� l� �T�,��c�-[�{��<��Y���"{�:7���w2�a�}�~uɌD*�2Т�+G��k�
����CSnX:��l�'�r'��I6�Fh�-��zzZ
Y
,�<@��Е��F�=�k<~C�29��L8?R����[�uP,l�=���G&�8�� ��I���ٸ&�.�¥�7�u�|
�$;�[&�^ʃth�ag	�>2�Q��O_�
"F,��l�n�7 0��;f��g��蓚΂�A�|g�}��X91<֓���`�ѧG$"�s����T��	��̋�?o^�� B!���;��7���i��t}�D�y>�/�MZ�	�����u^E�@Ы�nA���oO�0g^����'�L)3T0�K"��^hg��JV�����f�G���v1�>�b��Bh#�ټ�ZD���4v����i�5�C�LE�K"�7�pcq��Z*v$�p��:��&t��˜��ٝ֏�qQ�qH��C)YD�1o���I����'�+��g��/a06�᯽�i�{r�O D��Æ���f�5�U�u0���K�#vΤv�#:&��/+�NX~����5?)��u�^�?���B���?3��2����S���Lg��+L��$C��b��RQ-���G��b�̅
�����}�"�g" ���oy&�G"���wyvX��f�@ͅ��3򪂒�W���@:�lk���8��e���kM��z�-��J��(G�k�oYЎ����}����Q�{�Y��0��"F��/J�(Nr�Gåf�L���M~�^�Q�!~"��'��l�'���+ܞ��	dz'ĉp��M�^:s:WV�n����:߮a��I�qģW77�k�AL�'WЈ�]<�5/�V�Q�v�h���u(�_�����n^�:���=�� �\S�5
�$f<6')b1���=m/0Q�9����wTb��j���Ր�y�e���J�iTH��y��Qc�sPĘP�������;��Zhe�h�7����K"ߴn���
>IA�k�O�:�1٦1��,� �2���,0jĽ� +�'���l`&��Ax�!�$ Y/�" Z�2p ����Iø��~�b��B|�E����#�2� ���f%�L�+n�o��N�w �	ǻ������{5�}�0�9`�2�9?̦x�Q�C/�Q��u����%b,�O�&�H]w>�\�Ŀ�2����$�e��@;��KJ���H��7������vü���H
���)���
g��l���8c�����ІΪ@9OA�)(�l�͘4M{Q4b�u�G|Z���&�U)*4�� [�s��s�T��لW�]�E�E���y*�5�f���um3���#��"cַi�.o��Kg���+�@kC�z*7�J,o[�|P��/�o���iλ�d�$=�wte��Bf�����E�L��ã��+/m��/�#��[�q�jgGZ*�i�0;NZ��5V��;���܁���ѱ��#��1��'����V
L�Ke��kH)@��#��9�4��"�0��	�C�T �����%��ky/�)�ХX�\g:ˢ�$;ҕ / ���?׳�A>z�`섦��ZNW��<'�(���c8�ެƕInM#��,|a�K-�ż��^����SU��Q�t@�.�L��L����⵩��{Ȃ�����)�9��<.�2�L;�z]�&<�Ւ�e�F�A���#�����Hܾ'&~y
�6 _�Z<M�h�1I��L����o�D(������s9�l���9jy"�H-�f.j��K: '�Z_�3���q_���<��Оt���"�'�!�+��b8��7���s�ZA�I.
��v�3����@'�C+�ש�G�����P���/݃�V^���I�]o� �1ro�L���m����}��j%���HhY>a;!	��Ǥ	�GUt]hQ����r�O��&Qۘ�gJ(pm�#D��$Bs�W���z��`�g��7߄��.��^���
��U���s:xnd�./ʹ�Ϝr���K�$�g`���d]	QX�%:���@scڵ�	՞��Q_��h� �����C���?5&��F�?%�K��"tJ3.�a8�.���F-x~�{�b��do�Do�Uֳ-��]��Zd�r������MN����5e3��Ҧ[?S����E8�_z7��l��K͎�L�j��SK5�5���1�����}'��Q�p�E$���d����t�V�к��e��^[y���	5�e�SA@��3����%�����[ѵ����n��9�<�]���&��-��0-u�$���v����}a�1xY~��]H��!d]q{.¼�V�3��&j%CaS1�R���M���YK��r�ɔN�����N��ɇ�geI����V[��[Pu�z<�#KD�x��/�����r��Zk5�uV�險�k.kS� ����1�+�ձ��%ߢ(os�P�DI�5�p�|�pU
>,��1����r荚���m�R�.i�J����b�Оoz�-�CI�����q�7�����_�Ċ+�S�ʒ�o��Q}�7�����xto��?��
�vn�rӊ�g��z� EvX�/���!V� �6,:�Z�ku��-̤ U�vQ�_�Olyqp���m�p4�/�H!�YJ�
����t�%�ьx�ow�^�X�I>�'i��*��8�O�y�S�¨�K솜`;��Ձ-�L�SՁ���c�t�xn�ԙ�i^lb<X1�F�,y� �F��"B�ߋ�O0��[\Q�C.T��;"i>{w%X�<�1��X�*�N��6��=pj�|S�3��BN�YΙ�6�M�/۔�f´^y7����,9�.�ؑ1���NmX0� ��mJGl�I�T��Y��W����Nz�Ҵ��-IOrI/�O�q�_��.��QYN�q�Gq��>N���!����T�U" �)�-O$�u��Y�l�r�w�|���gq�Ψ�������9:}4�`�@��qؿdZBXk�&�N���D�7�	>#&�B��{-��n�Q�T���0䴛�� �C���X�̞��*���3N���� ��2��i5�V�d�h�O����~�?#o4�҉��oh)���LhJ8S��%��?��ͨ�uw���.�_�I�@�����QA�N�x�D�{�ī�[�U�����Ѽ[���El�G��� �
�)Q��U�Cq̰��|_��<+�L�_{z(u���Kl�`��˝�)ܺZ赬�Z`�{'=�/1U���_4�KJ)�������)x҅t�����hUTp������Bu}߮�sѝ_��~ ���<��dX�-����&(�><E-+�T~v0��ϭw��>�<:a���#K�1��WʓM�\u���A�'��T��m�k�I@��Q�m�'&��p\t2E��6��s��4͕LY�(����F���VZ�.:�7<��o|��XlxVHYEB    fa00    10c0@�ᵐX5e��=��Ȋ����ǈGFNϹ�E�*v�m>��ɘ��W��ż�xu[BS��V�����K�e���1NKu�y��8�C��,�aU��}����+��e���Z�p�n-�3ڭb
vZ���@�*
x#��0�p�w��HӜ1�Y�g���F���9�	�0�� /�=�0������weW�y�0q�r���<5�b��9ʚ8�۞&�`.
ӵe�����Y-ޟ���ի��5X'�8���9�Е鰮G=fk���A�$��Q)X��;S'9�w��\]r��i\��������vI^nG�_��%�W!.���Y�T�j��T�NDw��1����s�����j�w��a��{-*���dCO�=ь=�=8[Ο2��XC�`��5P��9L%:2�?EI�O%$������&u1�)�*�q����N,�S1�Yt�n�ٛ�;$�\m�i���&�4=�qX�4�D,�B��`^�]%%J�29�����T�~�}%��JN��Pz���y��An>k��q�*�{S�L���;�ߡ�d�����*��h׵��C%K���AD�a�\��\PJ�垽�Я�����N��6/����T��3"z#=�@L�vR�|�F~W�b\�W�a�؟�K����I%�lb��4$�o�)u���^��~���%q_�S3J�(_m�<�J����� �:�<R�x�51����#QJ4�Ո*^g �F��I�VG�&�a��d�Jw1I��=:�=�l��:μ�=�ʍ�����CL&�۟w���ad�)2�L��F���x�?B�ʸV�${�,�F��y���K�T#���ة�L�/��c,K��s��6����`�S��i*���`��'�����
,�8���	��`�oq^��a��׎4�G����&��	��{���B^������/qA���ҭ����I܆�#֞Ip��,�q##��̵�!���q�>�r������Uwc���8� 	�v�a�j\��[��J36���6dl<ι�$m*�C����g�ና|'2Ɠ�]6-A#�w��;2Sc}o���YlK����=���d�uL~�A'�fp֧�Fa�I�_�T��Z�s)�
F�<�_�a�����1��=�m<�S|̣2��7��o�}�OG���up��"?x�U<��9b%%}����O��j��.b����M�>�E�B/��KO>$���a4t�սfz��iLS��2�����D�hk��Pa�q�gv7�؞Z	)�vqE~9qAP��]��R�^��}#��vS��U��a��A_��͢����O7M� $�x�1߳Օ<�i}2,���C�*��-��+ox� ��>�"�$/��sr�{Ez8�iU��>�mJ]8���`��m�PO��Ex�'}�M"��P�Eb�aϗE�IaA��ǘ�Τ�D�gS�����#�)�둓�.ƫ,��'�/����~mk~���r�OJ��o�����E�����L<��Z�%̂�He6�%�WA�N['�؄��S�B�ۣ�.l!S����P�Y��N�����wv���x�[5!ĠNo�z�Vâ��>Ĕ�x+�b��5����,�&�8"�Do$��C�5�>�9֚�7^V~�B]u�����z`7ی�I��Z͇�u����]��^<)�t+��uØ�1#�4_�v�oʀ���͟���4��%24���AZu*8������w��"mC�ur�Ʒv/�@$c��m��e���cm��؛]d�~��9ls�'3>�_-+���emk99Vh��O������Ԯ���X���	f��Z�K��S��j�[eԡ"N�&�ܬF�n1��F�,=z��f�Fs}���Zً&�:���>����z�b#i�^Ll��kJ8��x	����LpX������f<$]Y��xeu��fHt�o<��.П�����Ns���E{�p���H"�˝�!��驎�ft^e��\���TKXn�;��P��5�z��*���xzN"\��(�Ǎ��q��?zY90	\+m$Ë��(HN~YDZ.�e'f����ě橂�d���}�y�a��M 2�'���ǝ=���������Ʋ�lD��^�x
bra��e��r�X7��({�iד��+��ӄ�M�1�r�'�*�=��������3����~�8�C)u�]A>�Ƒ�gOp����S,&�S��2JM��5��Ȭ C�ć��j�D�@hc�5'��@NM����{����xd�~�t�f4%~$&�h0��w�m�.J��8���Ҹ�5�J�`�%��7 ���w�?aA�q̺��K��3[]��B�.���T6@w]$e�Т�ֵ?�*���F�ǜ����#���	�ά�`�GSa{l�2BTM�?���8�N�3L���3���n�����['�����<� }.�B�!�����~�7O� ��ڠ�=[�Ϥ���_�|3R|EP,��~j-�˂�syB>U���J��en��K��9�Ah��6[+E!{?�}t���~X-^s�����G�W}�I3#��c��P���� �2���ɡ�tÒ���R��!f�ff�SH�U�����?�wLĸ�2��x��~Zt	B�oP��JAxPv�1�$�?���2�!���(��� B�����vRڑh/Y�sK�*m!�xO�:�x��_���O�7#�nN��m�o&�z(LУY��;��q����
5�Q�:�}�֡���A'�%��<i��ݒ��.���&��_�}0�?��w��m|��H���R�]&ı�7�\� �Ժ�ƻ��H���֡�v�Fh��{�.FV�����P��g0���HQ�Ǭ�L\0/�\���C��dk+#��.�d_�m��4���k�$�t`<�+��g�9��Dx���X�+|_[��� ������]B�}(�k�e��������Y�C�U=$ `-/T�i���1�G-4�q���+v�u����`�kBZE�5��|�:Ĵ��{f�������3JY�o�~�'=:������a��aV�J�O�c�O7���ә�t��b�����氍��� �z���u�(�l��b��uj���٬�=���^!L	��e�҅I0�`��:l�m����3؋2J#��W �
n�I\��b��5Z\5�?��D�
e�-K��;�O+/%�N��nL�"���b�;ҕ'�f�����G�ӯ��3"���TS���F2BvQFH	�_q����]�Ӝ�h�����5�VF?Q��a0�u�
��#'���* �? LI��D9"�ߡ��r�����wNH������䥾��"$>�������|=�>p�V�W v�Y�{����h�Yv}�T�'y�!3LO~k�y��} ͸;��a��Ր�+Kk�)�3��t�Q�T�)�`ذ����	�au�;�%涩��� ��w�n�<&�«�5L��|WkM�K�k`Z�ш�B8�t�O��堁�4�[�16 ��ID-]�+֖�����L�TY~��(���V
�V���Q��2Gu�1�v�V���h�͒hɞ�)ɤ�l����z�	�?�Y����`lwve5l}]�LM����R�r��OzY��W���7d"p�p�|?���֝P�u'Gj)�b,�m�����w��� W�ͫ���5V����������kv��MH��0���i�o�Y�>��Z�$�u�ƣ�^a�U(�����5�j��RZoy���K�-��~�ҺW���W�Ca���Oú<����8TX�"�3����C�(Ҿs ���4l�'�����+��!$L`P����j��E�*l�Q9ؕv��9��� }5@�4�c�I�"����H�,.P!��l�*����ε��n�<>ƶ�: ���L�p-~:a��VX<2`V�	���Up�"Ш�/�C�ҷ#3SCO{��2�<�1�Cӆ��A�DvA�\5�4����鬆4�"�&���>|rZ�@���^J9��D�N9��z��3U���c	jo�r��=�T�v��.rJ��큀�3V̬���!��H:��m&��ANµ�J�N��-� DN�.Y�:dz
��*�*}b4)��o}L�eX�8��H؜쬳�f~2�W�k�΄��J�K�u�L���}�9�g�̇��	ȳ8:��}�oE���w������>�	,E���Y@�]e@|/~�[m��gF'd���;��(����c�:i��8XlxVHYEB    fa00    1140�6��[���b�$�T����ӛ���PjB*������a�Z5���:�T;��k�+���Q��&�,
*����ኵ}�Վ��D��n����8�L'�����l"6Ι�	�����)����t����T�f���݆qIo^~rȽO�����9��yV��mRs�ڔa�����J-O�\��+���mӀn����n��E���R����]��#�dz�+���b^I���n�������|'��!)9�<Ww�����_��IT>�����t���*WfvL��@��vXQJ�B.q|����c˂A���Bm}d�/ѰQv����v�X��E��F�D��Y2��t9�R?B��K�ˢ�^�����W ̅��"�w�dI�t��%�Qs&1I�_��9>��x\�9$���DWz�#fb6�e!� V /����DքH��]�|�� ��n�a΅P���T5L=���"�l�-oȜ��",�HR�<���?9\������Y�u�O^I'7i<Wj�X��&�s�1�D��/rL��k����>n��,e<����z^ӄsv�Hg�&~T+�s(i< <��D,�˵������1i�EY� �� ���1o��/������pw�@#9-~�F��@`$�ǯ#|�UÛ�8��U�@���NZt;I��u��(@��Z��D����[a`�gX� ���n0g��i��E�UC1�\�+���_������B��
m�V�\F�䧩bG�L-�E�"���K�.�B��=%]��?.�<W5`�jۘ8v]Z�+�U(��$��|����^���Jg�s�(�՛1^ �PS��.�n+�����B5�l�6���sW?�q6�u&�MMI0`c�n�ZHH��s�Z�O���^L T	9���#����t��ϑ���(�w:?�B��w}?+�L�Zx�F���[�O���{��!Pd��Mjc���,h�(�ֵ���4��IX��z�B8ѕb7�{S=q���^���Z�5ݯ�����(�0�?s�=ƥz�h
cҎ�3����ܻ"�����g����[NaAcu*�-Z^!����/�Twt�[���C:�p��	{�q�\X�1Prsϰ4q���[	���ta+�{���n���+�F��@��(�BhU�ol�/��qւD�5���է@�{5�	�H=���\Xe��6��a�Z ����.l�����@�`�^w'�AR����"���Pԛ�ě�+�:G�y����+�P�;퟽���O��	k""�B�Q(��%���F���Ze�=��P���s�	��m�E9��֎�R�
�m�;O�J:k�dG�CÅ�q��&����V���i4VRR*Og!Ӓ�DS	cd�V9ͱU�L���x'�eS�D�1�jc��{��MG��GW�S��
�[�T��N�۹�ƿ��hFs��Z8�թnVE�e��Qo2ʹ�p�O�0#n�BҫY������|���F���`DX�o!���*�\�ȕ�Œn%d�u��P��CR�YE��\�v9���g��K�Zpo�����M^e�%�ʻ�+e���Q���}��������L�φ�@����ΰ��n��~4�ė`A��l̥�L���R��g�̢7��A�xᲥ�>�=RF���q���C�q-@!h�?�fu!d7�o��ŏ~YF�ٯ�C~����Ξe�V���(@<�2q��P9��eY�� �?(�K��d�1a�Q���0�� EP���/H�I�ʪ�9�H"���y q�@f�z����P@��+�!�Ġ����0Oe���~���_��|����=�D�k ����,��sb�'��n�,f ƥ�k���o��:�
�ėr�d�6M���l�Snl�Z<]�=�/r�c(�ٰL��B58^
\�^fK��/�K��J���ؔobP�蠁p 
�9.�;�6���A��]��%G����R]���&�0����� c5z4r���o�q�w`&Y��(Z���(i�֝3��W�z�K�����E{�7ί��>g��Sj�y�P�;��k34|~枇���Ky��O맯Imy�oNOl풮F0��4�:(1n�iʜ�u�"�����i����� xiR7��~L����r#^���[���o�h���-y^�0|+�9�y�z>׷�G�@��ۮ�d�2���C5�3Wk}1V��l�ۨ��t+$.{�A�p��s�,�ҟ�3�7Mi���D+}o'W8�
N��ױܬڔ��#����\Y�W�Q��:��,�~��C3��%e2���.f�uiF^�Y7ʆ8���Ì
��}�i�{�w�[����_)�Av�����I�`� �yu(�P�[�v%�I<dɦ���M��o1�O��ciF�t�9���%���Z6�������]v,� ��� �?�Oa�#��#m���������yg*�G����#l�\Z_0�S���5ـ���4��]��֎���=�s|%��7>/�!�^Ņ 5�7��(�2p�Юm��n��.Y>� ����G�	��VL��]E�K�+$�Ҋ��Oj��3�c a�c�s�9,���TB�R��^��Y��B�
�ݏ�߃�nx��suo�G�c��1�/!�5���|�>z|���%W����-��d0+��SE�ht��Z�MF���s��ZEz.�%�Y8$���%�UE��>>���͗�K�)$@}7�c�H/*-���a!�\H�E��a�J�@����Ng%���t��I*��"$2q<�}E#�D��0v�k}
q���l��E�_��سK�ħ�uq��O��A0�x��I���6͉;�<�K�l��͕����xB����.���k� �O����'^2��#s����R�ǅ[,�8����k�9bʝ���{(�i��lAd���3	Q�X�%���8ӧ|ҚGeSۂ9k|`<�U������i�����6��Uh��HnJ  5y�;z��b_ꃡqKz���Ӳ��I` -�\"E�&JA9����&��_h��(�`�
�	G�CsxƳ� ���L�ז�,���I"����o
�;��W�V������؄��D��*�u��1<*���ŕ��YkI���7:�[Q��Gp�)�+G��F�z�`v�΃;��]]MnJ�n"��[�cF���շƵ���8�܄�:��dɢ|�T�N�(?��F�����rM>��݆/�� �r�܂UIB����O������/��eЋd�*D����_��y�x�\wO�!��S��v�T30H� �#��a��Nu���D���ڨX�.;1�=լ-	���� S�M
u�#v���h�z;;�Se�+Onf�BpSdSS���#6��9)(��������ʤWؖ�'D�l�
�%i4(������:�p�"eYf�)a�������As3ᚦ�!M��T�ע��\��5����;�v��/;��#k��yP����@�?+&Kr�Ĉ哪�����Z�`A/X5v�D&�K��W�5�ܦPX���V.���ւ]l�=\�@��|� ���S"��.���=D�oٷ�D�Y�Th;��H�6��V�co��PS��<'9�:�գc=��|Z���Z��@�D�M)�_i\S/��M�W�~vb�YR�n|2�CG�v�*L��zP���6YJ�h���à3e80����D13����c/��]�.�V�!��S\�ځ�>�A��آ+>���iōA�JJ/�_t|&xW���N�����~t[�Z�)�d����MU)
��x��g���\l/V�Y�pG���C?��DL�g ��1P�� �(P�7�$77�J��Z�I��^*�%�|������P��K��� ���X�R�O`��A��/G�yYI�4���%���<�)���n�`P��l�g�R���6;�t����"��/y{x�$�����o�	;���H�I#�Ze�:"�0��-u������QU��9�< ��>-\&j�a�����*�*��G<F�N�����ba'��(E%�q����,�N�J�Ďă���D�b�{%*�� &�H l�|5O��<0p��!�����>`�7Wa<�1�Pa�ZKE�_8=O���k�y�����歜�c,������}`���2�$��"ڶ��C,ٔ�r5�+<��5.�YL &ú�i?�[�s4�@��:M�5�$�ՊBI���*h�����B� �J�^�2�=W)��uS�3��FH[aխ��c̱[ND���wf��т��-~�h�1"�V�R�IG���) ��EQ��
�!�_�oBqi��^a��B�{�� ��W��r~�x7	���+ܫ�.�䙋߇}�f�
?��XlxVHYEB    fa00    12e0�k�o�K��;=����yp���0���y3#Z9�9'��zߪS��Ȃ�4�
���'��hM�����y�'��_�L����(9P���]4��EfZ-r��q�Ez�)��$�Dt<�aw2��Ӑ��<"Ê��a񎥏��v'.B �?�E�v�4J-p=ڹ�ོ儝��knV���C?���@�
��L�{va)�6�������Ӿ�#I�ğL�����]�B]@F��DX�櫫i���ng�F<�~��gq��.�� ]w5��#�I�栎�?��q��g<����1f!�7���>!)؊#��Ġ��*����T��BӍ��(��I��Ȭ��*���K����h��jn��AS�/n�Wi�Β	;�Ŏ:5L�kd���2|'�e�5:��%�"8���Z_{��Z9�QCڞDI��O���D<�:?���9뿘0�Rc���I�ر��eZ|�k�Ϝ�7�)cjG�ز���Y���������Y^�a�1l<*�1��2�<�v*�|�H�8jQcL��L⥞�S�&l�m�D?7�-�r���o}I�H3�,������{K ��(�10 
t�ֵ`��%OTƼe_۩�ӂ�,�ѵ�'�)�����'�F[���L��_Y�8[s��R�m�.�-g9)qLP�xR�1G~��n�ٵ��F�s$��bL�:�����F(�v��+�����;�6��4�h�A��Ӹ k��@W��PhS�Z }-e�󺫑z�wAQ5��*�t�W�ɪ�@������RK�W{�B���M�׷�)E���'h�>���t4Ɓ"\4��� d��j����`Bt�A]q������DQ�Ӱt�Z��q�R]k-[Kͭȗ&6U���ˍ�7c�~��2}:�H!SRn	�.��bH(�P�O%���_��eè���$��%�u�������L�X�)��N[d����\����Xr*�-Nc%�i�/a.E��1\ܳ���g��r���,�7F�K7�co:'ݲ5P
fB�-�M�R-��}J�F�{hm:�H_�˪��������'0fE�2x'�@�Le�oS.6H��ZR�����-�y�\�vD���eV�s(K3��������Ɍ]r.��-���M���0꘰�v|��c���b�*s��y�n>���}��I��	�9�[��g�8?�4���
B
P.�|%C�s%٬a�"
��g"K`px�5����9�KO�eeQY��J�s���S�,���6�:����2�y���c�H��BN��Q->�~'iL�SR*X�k�,Z�H[Q����˳d@�Q�U�'�YY�9��ǃ��>H�j��I:dK�+�^���{oU0�@y���"3�R��@�Y+}!�n�Dg�K�?m���!>���2i%��-=�y�0��T�qЭ��f��P��xஐ����X��Fbr��1M �У}%l�i�Qw�/����
jr��(�bp��)վ��	�ҸyF������e�Lhaa�3�g2eG<[T:�	>Qax��oA�"�y�k����W����:.B�����R]6x;����Z�wQ���Ihჼ��L̂��R�(�j�#�J��(\<�Ǽ*�ܽ�8&g���4r4ؙO��qb:�ra�4���1��7"�b!#�?AO}��#����K�A��䍉�Y���㤺��x`(уY�x�
�2��>�`�����>C �D������m�o�#��ԡNM������}:�i��L�1��Ȍ���Z�.�9RŰ��h"��F�m�����S���,�w����&j�\��P�OыI�&��s*�;Up�-�A�moF(Q�Y(#2�A�_s�����Wyo�?x����e�O��;#g�^���+�-}DBPރ6��Ы�*�=��VL�t�e�>ī1��ǧ�0��p��MN}׈X����k��1i`ʩ�,��1,1V�x��O���볭�J0�H_�M?]�LD���2��̊�E�7�a*��!�m�o�c�+����Ŭ���w�����H����4��Fǀ(��`{�1Q���cBڥ�� ��3������1̘��/�BYC���<g�#-8��{Ж�A#3Ĳ?N�F�K[�{���#X�mц����#8c�ؾX��uh�s�[c�Y1Z�y�&�g�8$>h�.����]�ޅ�j��,s&d$�@g��� ���	9��St�����D�2Z�L&L=����|�]
ҋ���||��c'��-��3
r�0b��o7�"��i{�� ��k��V��4����Y�)�@��U�ZFC�oB@O�Y:��vƎ]s�i����:�7��Y�
�H&4�l�)¤�xv
ԁS&���}��`h����Ql�����{D�*ۜ�ɽvL!������Y�c�y�Ԗ��cg���: E?��m]��11����F-��ܤ��%#��~��Zb�OS�C��G/�B�5=�4��@�����R8k�"����ߘ^e�3S��;H�ĦDLr����^���7D(&�3L�('��a�ӧ�m��bI�4m�a*�"�$�x'�����?ͪxK����c-�/j�Wؓ���o�潴|�dMo��1Ko�@���D@c2+��=vR�5�:~��k ���&P���]�ݽ&U���L�/�",�$5�j�U55#�_h�z0��)Bgg�k�U�F����2v��P�5WO�e�J#H|�Y�J�L����[P�>�����<�}����K�ŭ1��Gm�*5���ep�!�$z�	�M��A�s����)�S<b�B��1p2�Woa@��G���Q	��F�5:�9��;�x���s_��~HYU>�F�'�ؑT/��1�q�Qb�T�H^F�L�s#�~�0��q|"�*2r�=�B����&������e�7��)�\�C���\`��T�E��~�b���Q��V���[�6�������@>u�?U�o����b'��҆��V��o��3�Gnm���fb��j-.-Z%'h^c���]E��a���u݀�
��o똼[l�/���+� #`<d�nI�25��(�|c_n�;�pG��1�l����C�L �V��QT���IJܼbu9���y���?eP���Če+`��Q��Ђ�N���5��ԅT/\�v"X��b�����F\ޔ�.o�{o$��}�Dyz���:���� ��o���J3D�f7�%���0t4:c�J��?�MB����Њ�p�r�]��օqA��2�s=�G���bav܂����K.��c=˺��TF���pXuL�]!������k
�ε� �6ͅ�J�K�e��Ч�R(���&A��<��?�c�(����#?�:/;����^�T�$�`z9G5��b�N&�t:d�^��P��\�����X]	��}cj}��ɢ�	Xڻ��wȮ����8U�R��������7fOz1�Vv���󒟩����b�+(8�v��3v��}�+�̏Z�4�
_}�H��	�\���u�	2���ڻS�Xb�,;�{�L���n	��:�@�2��2���C�@USkr��$��۱�ũö��1L��#�O�Olf��8B�}�fPR:B�Q�K�Y�<6� >��)3�L�e�c'���w�]r��^(���#6+��G�T�'���7NZ��X-M���0'��IF���[�S�zj$G뻛��턶f9d3)"�p�\�:�����

�3��0
���jbxg]�e=W�x�Y��YR��Ti��+��d�3T�Xp\|y���~7�U�8����e�_�{/��(f�r�q0�Tu�G� p+lאc�j�B�Uo�H;�l$홬A9����4������1�� ��_����b1	� ���oI�&N�����k�fM�I��<4[oSG6PiXGpGt�:��*���ϲM:��1!F��_�a:�Oa��D�:����Lu��k����t�N�عE��xݐ�m�vM�������(����ۅ���w�`�<*��u���M��V���dd������f�E�i����ܒ��z�5B:oű'o���ޭ���	4N���Ί����/�Pk�Yfy��d�Kt.Bo��d�8Ʋ��`ȤD�-�|�P44c+�T���V~�yeWm�T���j�Q��p�}����L��׫0������嫊&M�I��b(n��ȋ�{��عk�U�z&���^��ǤTU��D� ��S��I���!�+p�Ч�SG����M=Ĳ�e��=��$���Yзn4s��9��/.w����MF���l��=�M��+G��x��~�j��B����Jm�CE�k�:� ���ef�����S)H�O�Q҆��><��N�m��1���]7mdUA��!�D�M����A��v�ƙ'
�P �R%����DW3l�� rj���%���:�:�~�OƬ*1&�T\&Lo����-E�	����|�{f#����pc�S���V]]o,=�rI1�$�'a�Ȳ��_�PUD�? �slvO���*U��bl�m@U�.�1��Bk1S���S!O��UpV�aິ���d�3C�Jh/v������62b�r�H?-�bJA(�i�k�.~ax|� ֕�kE����~"�璖����2�e�NE�|��j�@��.�8�a5��d��n��I.�\���g���9���/��*@��w���6��=n�9��\�ϐ8�
��H�D���Q;&4���v6wcd���d�.y���0���'X��ݣʁ���Ђs���=�7�-0�=�>�w�C��}�XlxVHYEB    fa00     f50#���S�ҶɺJ�kW�l�}�9`L����9�ad�ɟ\y����� �H|�i����G��U�b"��ҽ�����6�Fխ�ڸ�5uW	������d��ߓ7V�;$��<����J���/7VY:�0�Ώ�g�?�rh,e&�n��q'�u7m�۸�4���.=_.��ص�΂d�Hsw��w0�ߦ�����93����{U���n��4F&�����.���D u��!^ߍI� �8Z���$����&,��YK�@'�Co��X�}��u�{�$��P��a߭_{��Zp�z{ܕ=N�2�������n°�������GR*����.¸�)�O8��=e���(ZZ�+4V"�����pôv{;������<�8�G��ҼM��}w�l�$PB�<0��g,q�l.����� �\?�:��k���8w���,">�Tz�oS�s�(�P4B����Pe����gG�;2�Q}���U0��Ro8��� ډ��cOA�.�L#���"3��,�L=�e��/����Ô����3�/�.f��/4LlB�T�.V*I�����G��X~�q��;��'�k�E���,R��E����.%�&j^��0������>�Ů��s�����ع���`J��V���R:��/��Y���}��&Jj��>K��n���8X0��!Ifd�W0���b= Z�k�<�s�~j��Xk��L��;����w=��&���H��&���
eZ19.�oZ�f88��兊M%�ҥ����i{� �)�i+�'��Mx&2��q��_��_�YuwB����H�,�s([���@�]��f6tW&�̨�.R=�pG%��� $�;�����T\\�Go��� _��l�
� \�&'{��J&���9���<�Յ��z�;��AR�Pq��
���a�j����s�Z������sy���մ�_"{� ��0>�"G�3Y�(���`&�ʪ��a�L�t�+U�_�h����!$��TZ޲��I7I��0I"^J(�偩��4m��;!�'�&�\��[�R&�+ݣ��5�Y���^�^�4�K[ރPޤ��;YɂCGg��wR�c�}
�l0 Q��-��M�#2�}Q���;D]�sKؚ�9a��;e�s�X$���1�v���OR�|8�s0F�Mj�^?�r�b�^�.� �tJ6�4L�@R��h�h~�T� #Z�WL������܏d������
xR��*�\�?���De�1���X����� L3L�@	5Q*L�(8����w�t|n��{�z�L��N��5h�,��Ks���2�ŝx�#�~���&���y�CA�9{��ӗ��jY��4E��_�x*hkr�:��.�]G[Jt�J�C�H�������c��GA�W�R��H^U�+�yaII��y���.�ǁ��me���>� �Vx�I�� ��]�Z��ثwk�|�A��c(�������*��0zo�c��#,[�C�C̸�{��o��ř��,բФ?�{��a���I�U���YZ��Q����^��s���f�G��������U�*>����}'l�5������5����kSk~`.�ك|c8��퀬34����G�_t�3ǟmc��f�~�9�lS<�2Ȁ�s���Q`��$�>�-)���G��^�$�d��G��Os''�/����QUJ$�8�ۨ�ms=BA�F�>?�Ti���r��^����� $7�>���P,Y֌=64(V�5�I<�;�(#s�s�KC(��kU��)�hT���&��
�=�t�t.�v�cR!	��%��X�tCĭ���p��Iw�CV��*���D�X��O���x�xw�hg�q�Q�H_	;
����SU&��8P���n�E���7�>�ҢZ�� ����_5�d#�Ywx�9�jQ��:YX�
PO/�1�/��Q�o�g�*��]�`���8"�	2v��{������V��ɏ:�.P�t����)hMɍG?��~��7w�� I�	���@����=/�oO�*���B��|�e�Ge-k@ �p�d� ��âk����t���Ƀ&�b[u�sܝ	(M�-p�;J����I��JR�;(���&�VE7�����Q������\^k0�"u:�Y���a�01�i�џ:�6�.��j,KJ��Ӝ�c�Pp�J��pn9ï�&�p�)GU�P	ۋ�����ibv3�ƈd��u���t�3R�J��2gdb������0.&l+M6r�k�o-D�T����$^);s@�e�.�L`6 �"9�֜�"�u�\�!�k>-�{jF�Bj��1{�нΝZ�zw�γ�%�Nۖ�>����%�e'�[�C����e�PL�.����ړ#+�s�V�"��,1����(R�t�o�}��r���?La;��o�p���P4��Y�1z�����C}э-�1��J�cf+0�g�"�1=C�Bj���=Gܦ�S�����s�?[7�@���|Z�61ZM�j��[̀�s�:1�g9Ak؂$,�냑=�R4N�mt4��6�����,:\���7�q�| ���-�܌�/�����3�T$���_���A��!�UD� �}��V�L4�]�w����ݘH��^��Y��̋÷5��㻵�}����+X�G����2�+"H�~�l���L�NWy��669���.j�L}�:V���Ә�兪�5ڡ��4h��x�1t��r� l�ݝ���L���d�:�x\G���x��#���R�j*�̋���b���4O��C׀�W_W*7J�G�m[���7U9Y��ُ�Z��z���bT������؞�}Ѳg1*�:�e����4���>�\6��!��JSMX�{�����P�r��.���9I��gۜ<7gҶ���F��h���H��S2M{.�"�g����ͽ�j�����:��5�%���,-��E�Ģ��\"N5Y�q��Sns��vS��'�P�D<Wk�Nm��n\O)ܓ4�o�)�")S���ڿ�>�Ԫ�b5�LG���W0H���3��!�YT�$��˛Wσ*J�@5�7������CY�h�!�%�-h���t��hKT~]]�Đ�����傦^Ѧݡ�";`��.u���3�Ҩk6u��5�H?C�)��o10	�\2�}��ԧ��	���NzL��t�C�9c��bƣ#��-xx���!	0i�Â�Oc�hf���h���)M�L�Iq���(�^�g]���e2�Id�-�5g��	w�v9k=��ϸXf...>A���w�}OO[!��$nS��iJ��Юsc->3j�{SQ��ۍ�b�)���q�g��I��@}!��bA=��e,��D���>�02_��(D]4�o�n2��&h���v>��d�c����$}b�#\N�w�~��m���4��[�I`��d��'���)�f����RZ���KB���>�_�[���������+���z�~I�b��s�(�sE�z�Q͇���;D����]��E3c�M.���Zv)"�Fa{߰����tpSeu�eн$��3�V���5�z�\h ��<'m��?p��:�=X������h��=�g%���+yec�Z'�A���^�'R��Q	�2`�gݹ��`���_�˲�-!Iwcdw%� �ߵĆlx���c�^$�&��4I�����XK����dQƎ�D�Y�/i�����pzyO�z��_����\���R�揼�ݗ�zY[ ԵSw�Q˳�
y�[��w���y���F�j�]	
�C��e����8RRK����H���P ��
I'��.O��I�bXlxVHYEB    7273     560�|�=�>o���6_��#���U��	Z�szZ�<,\-4I�`i��,䞅���X�`)��${�|��"d��䈁��Z�ح�	���F(��67%���[��Q�mi���g�� �"Ř���t��|/�7�����h�a�$�F�ɺ{6��
��=Hܧ٬#���N�����Il�bHY�0zP����X��8pyv>�p�h�[�{�8�f�z$����oe���M���acm7:���≈�sS�����툅p�5��D37�Eճ	-㱄���w�$�ʚ9r�X}��F�&_ʞ���q���1���[�DS^�+SN���9}UO{�'@��h��Z>�΃���ӎ/���!V/��[3_�X��҃�I�Z��=VE�}ҽj�󌸮��e�E��%�����|��;�"�6�mSm�E�eQ_� 
@�\
���j=�mE;�� z[����Jq�0��ۑ?I���I�`��6�	A��
�v�����4���`ʮyH�8���f
�aV�����Ǧx�3ӂ{�#�s�R�=���au|��qEQǅJ���r��[�X�M����yÄ<m�-P
���3�J�*�.�[6ŷnrua����]�8I��J�y�CI> E5�a����hj-�q�Lr�����\���Ȣa;4�a�����v��o�.�s:t���/�|>� �E�R�	��0���mvZ��{e�jA���³fze?k���o2E$����
'��LɈ����#ї�x\���(f�������a �l�y�N&O5�M8Ya&Ж���Hc�	
��*���ڵ�����6�Q��.��/b+Z��N#��7�G|�,��q8�kyK3w��v��w�3@��:z��;����v4��;D,BO�z�A���a�H�J�6�/>�B�6�0�2�p2�>J�Z܇��A�^�="��ޤκ�����__���������\�fo�ۻ�"r3;fRyףtu��`�:)�P���p=Hz��z�:_xa&������@��RдR��ż+��)�vD����u�K�BO�V4����:�4N�
���)�3�u��	-�n��Z��xS�%�q�\�%��� n���N|���Sx����KOβ9�s�]���]�a���B5�^
]�Ys���/c�\��(-,׻���#ӡ.Kz���Ā'
_Ti�+�k{�	o��b�S�]��C����W�u0˱Z$�[Fo��ݲ�m�岁�fH\�R�,F�t�s��A3�8B�5*����)���&SqF�ngG�F E@���ih@KaQ��Q��cU��d�>F��̊�[��6G�5��l���X�2��*r��m�
=%�ʹ��}��==Q["f�d�AG