XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������&�M��3\m���$�m ��'���m�����H��8���Q�4�pLSW��G�q�H���a�:�J͋�
:A6�^���V���>3�W��l�qo��6ܰ���ZOHR��t��L�'k����g�8�3����� �I������=@��h���y|{�u��r�]`)��(h���hE*�R*��C�8�^Q����Vఁw4�~��ƟL3O�c|b�"Y=7�xH�� #;�O�C/U�ɼ�{������/x�	Ų�z����m��V�ٸR�:���fT%� �f!�� �
Z[(�;I�Z�<?n��j��I�*���uj�愎�|d�q�S߿ A�>�:�	T��{
���6j��H[��]���r�4��Umb"+��^	��CD��0�/uQ��7E�#�?�;T��S���<��2����~cg�$X/�V��U8,R�-�͝_����&ςB^�]��֎Ǆ��d ���6gT�RX���Q��S��d~��B��ae$k���� �9f���'��e�/�CF�~�"��4e,f7	 V���>�H^ �#V(А�[h?��Il7Z�r�*4}�V�㠴#ϸo�v�%J�ڹ,�O�r�خ���^�{wL�l�c�� h~A6�H�	����uj�њ�>v)��3�~��{̤�-o�i5�*�4�aZ%����,��Fٚ�+?.�ʹ^��f�-m�<��t?��N����y+U�5��0��G�uiU�l'MXlxVHYEB    55a7     e50������4rR%����tZP�2F=}�N����_CNS���p�v�J^��O%��§�Ȟ��k�s���"��9��� ��� �;���.n�����n����Gm�V ��7Zy陂E3�s3�wL®FbD������&�
mѢ�jS<�w��/���"�_O�Ǚ�r`���V8���d
�w-�
G�D��R��-�4�"�Q��X�|^\�mo�w�[Ƈ�V6T�|Mw�V����%<{\����U�r��]5>|T�4L=�O�I�M�M�l>���
��7�������RV/|����Q�؋�#`��ڋ��)WL`�J�F�'��2�,�V�=h��f5~�]n�f��`�;�?��>~�B+���}@���=4`��߅=s蹮�ai:����R{�1T�A�����.��RU�Z��hsHaG���FXB��b��:��*zs��c}U%�ȮQW�W��{b�6!چ�����W��|Y���m��e>��/DS�a�	�ȑ8���|w0�ށ/�x�zߪ�H��~746,p����L�!O�9u������	?\�LTZ��4B �É�u�J��`�:Q�h�ʭ��S;_�>���o����7�]��<�VQK@��bO��Ў�ح��b(�ܬ|1�f�@��|����*��)�8�6�ƪA�P�\?�ś>��N3é352��}�����
 �w��gd��������\%B��
����gI�;PT���G`�K��Ɍ��a�=y���tn�P�^M��V謁���FJ����N�pX8�V��d��+���o�@DB�6��&>��,�������`%jf���wZ�j\���T�+ #����i���7��G0[��[I�n��y���-)&V�4�b�X���z��$�v�)��-�0��VY�'q�&r����K�q�$i��VT[Ԋؐ��.R�
R���q��jŭ�9����h��3�p�����9u�o[��:"52Oh�23Qn:~����"r��̶U��Ky-����>�o�j�Ȍ��Ҋ����6��R�b��eᵝ�h�%�n��5���ia\���*8�/k��EW��N���;�$�-$RM��[_� 9b� ��)�I��zX]�tUO��l�m��4�r^�����?�tg��Yt�[��R7���NH��1MyA,c"C^����:;��;��N��Ck�e&+�h�e���3��AoV�J�t_Wf���38�{�a_pt��s�є�$�!�J�>V�m���/����#gL��*Tז�D��oL���/��,�$e�(�O���W��$D�?�Hb�1�E��5O���5k�h7�5��jd���,��Զ����4|]1Z��&F
��~�1'�)��q�ؒ?~$��$����.�f\���C�g4z�5 ����VX��A�L&�"ٮ>Z�
�"X�D]&vO��r
��k��V&�:>��da��I�R��/�>'�� ���-����{a.C��O�U��Z��	��X������!�u XC����ƥc��N�m��f��w?k?���}��a�4fnݓ����Wq���z�����Q3��O:��$*^������/���s
�i[��h��G�F��k"�@*VTh?8�%D��cJ�2��u�з��R�m.aMHzǛ���YE�1 �R�+|������V�]S�\!��i>ևlf�4���1�M��J���5����y��p�����n(�QK�e*�\8��!2����"퇺�<��=#���	��d��e@۾+�	�2sQ�M'��￣`P|���C`����^�۫�t�U�pf�"0�]�����~�q�����wObK�n�l{Ys�K
EWB9	�����Zo�6���j��i��&W9�K���+�veؙ~�:������*�Z��;O^��z:�2�r��rJJ��,�W{���@<q8�Y{P����E�$Α*y�H<r�PL����5���~oԌ왵�]�u�׿�sI�,Lԓk@~�1eg`vY������b����e�c���2;�)Q�Cz��N&��:�֦�?�,o�+d�v�*\�@�0�سt��L!���ћh��r �Ʌ*
�S����M���F�A��jVA�Hc��+�{4%�јl����r����/n֬�6U�?g���,b�W4׽=���H�[�p�T1�n��'�to3Jͺk�RG0|L��z���'�p�~�`'/a:	��g��+@�ȥ�oӳ�y4-[%R9J�e�I	 ��_]Kht��_G�i���2ec��Q46��,�?8d�D�lv1��T��Y9S���w�`����� �(��
���n�S��Ͼ��FEd�S��듦�� ���#�I�߯��ͽ�=g�r��k-�P2�
�
�#�����<�k�w�E��<Թ!��%s��?&a���wh�k��9�#z�����\�)�S�&E1u����ip��bJ��;�"�@�Z�w˔�����s^�f�6��0��Ɖ�Z�G?�A�a�u���:�����b�1�w�F���sZa�΁*A,��Z�4 Ј��K��؇$�����p^�+͘ȪO$�l�~�v�.7ꌭJ�qڈ��5ix �/�x���V�������!X���W,��J9ecN��c�+�+��q�>,D�jCpoj�W
Zҋ�'k_՗��).�E����c��aS4@=�I7�}�1IQ���P�4�^ĚB����
�X���94/��-h�wҪ�x�bd�؆"ߟYM��,ɷ�'�Rgz�q��⳾��'��\;}|d�0ʝ5$��܊^�����C�-�Wah��x�������Fx����Rt<�$�ϳ&~�l6Y��Y�4킑��E�`�v�d����� I���YEK��I҅�,�	��@�ZݲU�����)�+�����Uu]$���k�fznC��IF�V�O^��������{����4�������E��,�I�C�0��ks�y�j�?1Ը��#�*(�oh	G��ta�>Ѡ+��q Rĕ8`ڿ���F;��J-��I�޲
��l�YR�`��r��H�&�7v Z��(W���X���yJ�̺������ޯ���0�2*�d�_総��,�Tr�p!��Z�]��{�J����Ĺ��"t_�c�s����y�?��;�m���	6�Ϯo1���S������2��En1L��ҽ�#�Wn����hM)�^��HM�ߢ�.�PJ���&'���#Z#M�I�0���Z@!ǹ@�l�3θ�����:�'��.ub;��aHtiP��Pj9��;����U#��Ne�gu"_-��I��^wL�����h}�ў0ڞ]�a�.�7���,�B>����������$�?`8iϬ��9:��` �2D2ށ=�TBk�݉)�m�������G���x��h{o>v���3�,-֙�Q�!�Ch�g}䠐Jo�L��j柟!����rn��۪��ي�lOyA�O�x�(畯����K�#ja�ɠ춛(�Z�8)����DN|��ДyY2�yN�4V����f���|?-Y0	���Z�h�4�kEG�b�HfH�')T?�