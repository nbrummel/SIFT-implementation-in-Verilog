XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������4�Z��G�I�ƍf��$����f!�Y5��i�p�Y�r;4�d��[3�ڧ΅�����Ws���Ja��╇�$�a�"Z�bX��	���{��:O�	�Fz�d�������N�i�£�G��"���`��w�R��{�OU��:�+�3����Y�=�@Xo"T����։D��ѽ�����C��Tb�F)�ָqYN{��T_��� i�ͽ��aw�z��3���11�\��"�i��c�c �,�zF��*�\xZ�WX�/y�l�%4�&ŧ�l���=�J|��k��;n���<p��*��¹y��{���
�t�_WL��N��F��ڄ:n���`˃����U+��g���6��汒i��c���ܥs��P��?1��i:=��c^���M����&q�����+^�-g���O����O@�|�F񆢍��L��*B�П��C%g��ퟅ�RO���q�l�\S&��-�1�֤�q����	���5��v��Y��mt��l����jЅO��M�V��:��k�+�i�]�����}��B� ��FJ����ߦ�C����LMd�Y���oַF�tSh˹�D�z@*cM"����)�l[��l&FAI�r�C�9��ע5W��k<0���GX�') �U���W3-�K�`�4�<�deUZ���ӂ��
w�CX�à��9�����Rp%��\���i4�a�|7>���?�(�Y���!$:9L�-��<4��^pGXlxVHYEB    5df6    1510?8<���*A�DN�Ï����c�vE���ݲvQ��tC��Y�W�|ļ� ���}@��TQc�`������|C�w���QD�R��{&��m�~̷���΅�`� ����쥞��):P�&B�M���C�laDAF��ٳ�<hI�C
q��BU6��tp8a4*
Iv�[��%w��$Ad�`d�RGE0'h�^���W$1i���Sy�|x��y<�1�M�Α䯒/��K�t�A�(Ȅ"�E��G�gE��0����}H�Y�B�t@jSZ-T�%�)�&"�x�8�Zo��q �ɜ�A��f�6���D�¨�J?���u�+>|���u/�'3ڣA&���ֽB{�%�NF��I���S���_�4X��f�]�T�z�Ѵ-/YgּhM�"�5ne������G�؊��AB4�@~ p:ވ e��"�MwAgؿ�o�<zd��ajW+��u)����>�G�-j��7ja:�R��d��$TtD �( ��3������O��yc�b�9�T��F��u�&���C6\�������R�l=�`C��T��R�\��՝<_(	U6��'u��8lz�`����a�!�jY-�Xi$׵��ԴB("��� ��L~�ѲY�@����`UuQ?hֲ&�jJ 4�UHRG@8AM�+���=O":m��j{�)�]���rN�.˒�Ê+�Շ�*js!�Q�y@C���۱�E7��$/�K�����36�&�,.O�#\�I'1��D_�L����#+��4l�8ғW�|f�3ѻg遢��,0:�r����W��	p	%����x�}(�:�3����N�xBR�ѣ�7�>��r٦�1�q�=��C�a���+��[W8�o���D�(jY�f���P��Tf�9y���$��VC���]�$��k�.�kmd�L�B��@�h�u,�+��hG�X��� ��-#)������ϳ�����=��y��H�p���`�P�~A�),�����f�<-������݂
��?��+6@�n�a�S�>G��h�1����o�).��ǆ}��؀��+�ǩX;��K	�{�-GJrX"������p��}�|�#ޅ�&�@�k�T���׵��?��A��0�n��y��X6��ߐ�:�ײ��
0���b�r&=�������c,Fu���π�l�|��;vx�`o[���07�ZF���eӋ`*D��Y��.o�%�\x��l����/�0�K�p�H7����R�Q�ݍ���2^*�2	��[n��,é���
�m��FX٭5�Z�g��"v���W.Y��sy廕&�n�ӀV�F^F��K� �]f�.�!�H�� 8��8��o��t��t,o7����C��4�Y�	��;Ȩ��F�?�?�[xO4ڕ�	���b3��2�� '�}�ն_��hZ��	c�.\%�4��hn�ս�)2�������}_�^�"�L����C���c��p�L��y8"�z�y�k��+����x^����U��j�K����%WL[\EL�\���F�����iS�t��Y��W|��K^Ѩ)��-��ni��>�Qȥ�c&І���0i�Y&��3t,���3������跬v���"}��v��q3l�����*�O��D���1����r�Vs��`P ^�6f�~/��_"�R����lB���P�5s�`/�Z0�7t�� ��(�遲��CH�D���'[�3��K}0VС�ρ޸(풭*���?�n䥫���]�	����&�����Ke�S�سivOƵ���k��\%?���WT��M�ۑO?�M�]4Iqc��z�,Olt!�%�����\v�zf�����.:��-��.�g�G���*��m���NJ�y)qRsޯ�����ůC5�������f���oA�o8����Q��k=�L
���)���j�何)hG���	V~ܥ5��P��
Ot�^Z@��x���}P�;���OC3a4�R��W��u��W�R�_YA/M�&���.+p'���%P�A*ٚ�V�6QH��'h��+5o+�p=)�19��?�~�U���>��i��U� �}���>V�5$v�ن���%�ê/��s��W �� 
�m���#䬮���I�/�������^LҬ���C���
�#�;	Ň�-���ܧ�Ҡ(���"Ta�ʩ���>��ך�fo�us�)�C��4M��K�$	u���,�ikhP���'L���A؃{�] ���%~WjP�	��P�-�M1Kp��?>Ǣ��'j^Տ|���uTGj��Y���ꛌ�/U��w��JFn�]Ƌ��d�n(L
��J��]�"J�П�yP���U�4v� a0�����n�uo8E�ƌ�}3��D���-n����,rf�Kes�:=%ϴ��'���8U�y�IfzCϵ�sF3�v�sB��I��5�e@���ƂU���o⟠�e+�j�1��}�CNPL��w���Mm���]�5׭GZ��;�f�ܳ[|���v�E�v�˪�!6#�5��Yz]as�uk��I��wذL)f�W����zmg@�3x,��+x���2_hk��zU|�*Iy%��(�n1z�H褵"ۜS�}���sѹ��]����xI�i�X�m����S<�`�k��Tx���l?�#��ַE��I���Vo� ���)�����s ������#J�?rT�!S��9N����!3�0���F{J�lDӾt��iI�����l_q�`���ҋ|�	���x}�$X��Qf~i ����6�-�;?���rԽ\��k��p��P��36��;��T��V�3 �ݖ�^*���&�2N^]���$(������LK�^zg`B��8�:3f}~���
~��	i:�2v��"R!Q�f�^n��5�8�	H���bf脞� :��S����>�s��������ޝ�?�/�M:�:#���/zҮP<h�C��#���	ˈ��#��y"�z枭��Z��+Ѫ������yN&��c��4����ҕԕ��t��U����:��J�A�O��OuoR𰘘Q���HCL1�E-��K��>�_�=9��Wu<
h������^�]�W��NSo�.l�yT[9I��%��*s�H�p��P�괙�>��׆�ϐ���~�}�������x��Y2���� nw~M�}�5��^��m���amtI)0M��`�{)����cm"(�0��k��J�7�8��J3�Om�;tQx�m#��K��oz`�BL�j
NT�z��F��F��`z/)8�è�ޝη�@}�mh�X�!"�B_��4�*o�O�f@�x�����㲥x�yI���ZٗD��A�|�ۭ�9鱎�����B4@�D��g�Ҁq��*��
.htar6��a�P�K �[�c���٠ߞ�>��G#�/^>���L$d�
��jj�p��o:���Z����^l��� o2nm�����k�P�k���K�4	ph�|����xb�-�j��@���4ŧ :A��'#yrͤ������!���� �æ:QA�nӥ��R�,�d�s~f�
!�$uw��M]�kN�����FNG�Fbu���Օfqs���@��Ybo+q����k�����!��N��h�����`�y� �&¤7>�a���^A@�K��ꤻ�E�C�yW�R"�N��v�qId�5{�P�g��&g�0���#��J����
$>��g�ЌK�dUFO��d
���8��^Q�h/�2�<�����Vڥ-��n^��ԓg�^�E�2�.�[B�3%4pA�������o���!���vLL����.�#���XBy�>��:h^� ���=�������g1�3@�ԑY�Q�N���c �,"��x��3�>�l��U��@G}-U��&���촌܆��,(����S����fzƹ3o�Q�ִKTD.� �׷����|�B�K�n��E�������c�k$-A�� �_I	蜧ňP�TT�w�*�c���yh��*X���W^�sQ�eYɈ^1%�q�~�@��|DO���f��Ъ!1��yK��n/�^}R��%w脎�?EP�o<&J�Ng� p�ы�iu�p�p��/U�Nw\Y)*���V�n�l���YEy�(�ǄP~�9]��Ǘ�q͗���������t�ā���I��wϢXWɜ�ql9�|�L��S:;sd�2�v�9�\�M��,��lT�'0_���]>kʙy��z�B��<:� �[ ���u>�6��_$�������=<�����^,�ꋱ�!��<����E�0�X�K��0�����N���+8[bm4�e�L_�A�i �}Ȼ�AwP��#�!Z�с�!J
�t%��E�y%��˵�����@�n�:�fQ	�_-�ڈ����T�NF�+�UThF�Q���Y�" ���D��Iv�;Vh�3����荎S$$��zU]o����"	��	��+K�HQ��p�":�̝:��᧐�h����ȠkH�"�4����,)���eđ��ҽ���gj�M���Xo���< �W^9�7@_�z�%��.ױ�Y� Xw�{%�q� ��A߯N}�xْ��$�.1.�wu�[}jgB���\ĵ_J�O��P0�d���u�z������ґٙ�O5ȵz7G�}k��;�M�h����t*�O��gj����p��Rro[��9�a��q�Mi���ܷ�.��]K������q���e�^$����T�!�Թu���1��弨�~"��_�`0���a)�hx���g�^�e-�ن79����bCL5+��	f�?�ׁTS�S�(|5�4�!3i�
�X��x��M2~�	X�Y��^����4�bL�WxRYLXs�4�?$�*i��V�˘w�)+8Ps�;��kI���g/�'��l �t!�F��=��L������۽ªd��yĂ����8uN�'�-�.:o�h̓z�'�uA7��R��z{=����=��d�	(|m���>0�@[����D��.0�߾fM����-��x��ɤ��|L�%P��4�ZV&��6/�z7} �N���R�9�������Q�g�3����u�خ�� Y��}|��D�i[�7!р��E�1+����I
�6l8	-��:�47�T�S/rHf�ưԧ6��۩2 G�kqP�T@q	����_���*���,sh���O��m���g���2J��Νb�G�\������~�e�"eF��4�E��Z��
���$� ]��_�-V�Z�+�Duxi�E���d,"���&��)c�{��<�v����BbИgQ9�o