XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���襬FCR1Q7����>Yj3�جj1�^��<wZ<��1�(�R7�%��/(��a�1�}�qԼ�ܙ텩o�gI�s��%}JGo]K�ʫ�
hgO7oqGמ	�
e����O��� ;�?�
Z���(~�A�Ф"�� ^9���C�+D�g�t<p�.��J�e��������r:���a�Ԡ��F���>��̼���2����H=Q2�Z)�p��+������\T�saN��ʋ�9�ĭ�
ϼ(s��ҵ�������%�U�/�"q=/���p��#	�X���B&��<_w��OY���\,�0R}&<�)���M���]p{��E�2�D(�{�nL���<O�JngZBpqse�ÅRX�h��RN�Еπ���\rkp<sC�q[Y�����^���ߖ$p��'��~�9��S뷤�R�˝�ǜ�%�rt�q�V�����4�^,@�7u�bŮ�\dd�Q�R~Fm�_�L��h��cM9C��=�u�i*Ձw��ܛ���	�۔��?�M�ه��ҰW"�7�q�*q�`�	���q����P���-tY��n%����C2��;	|9�ТFC�!�\�\�����t�b�C�K�I,��ݡpc	�6���*c�o|�uk�h�dujL�p>�X�E6P-��Z3d0x�z����$��b>r��r�N�WƄ�ľ� �{u�r��33{-�`f��uC[��)�s�Bd���눁=)��Wc�#�?�Q�c�@�{uM���e�qФXlxVHYEB    fa00    28d0&FF:�z8r(��ϖ���w�vo�35	`����Q��:��mơ���g10�xQ��$������Y?�M~#XV�0֋����B��/��G��4���m�;GȤ��ߘ�y� ���>�Y��ݝ�3�*�p��a9��(�M*�x�9k�\ġ��]7s����&�i�15j29#^��ˁ����܉ywZx84Xг5p/�`ؓ-k ��j���T�ȵFkP��@�x��(�/b_��<�_U
�D��0���$4V���;jA����'�^���Ce�Z.֝/�3Q�r�y� ���#�y�<͈3�6�ל�;	�qjϺ"�)����_�ϳX��I��R�}��xO?K�SN���k�M�y�:����d�y'M��5E����Ѧ�[j6��z�S���v�ڨ������Y{��Vq� ���|_E/l�LfF��H7��I��g�u���_�l�w�p�lQ�q9�w��ݟ�	��dVXo�Ն�oҫ��cl!��T �EZ�X2�]p|r����|��5�6�,�4�NKa|y�d�8���͵�p�����������:��������'Dίr��)/'>j�qRY`�!�X�I�vn$�%}���Bᛳ{F D�l=*���հ�U�9U��?P�`�sqd]nl���N���V_^�@�ݪRq��Ⱦ�^[+�T������mK>Ŀ�L�`�z�����ju%���R����n;�my����P�T(��7߃�b��(ch�f��6(駺�]ѹ�4=n�+`={��y��4�� �!l:��G�ǵ	�;��j�H�%���*�0KL��|]Z��|F/sYH3��>`Y�ڈj�ycĲ��*�:��9%��0�lp��g�G`P�!tN��5�-�q�M$�v��@]/�}�5��i��!͑ �2�ڿ0���91�L�1u!�B�5M)�J(�>6u�k��4
c�H��q`wy�By7���H���jwד�[�Z֜��������i�ɛ{%4���7TK.@�VLS:���wسe��k��*~�f!��WTp�o��6j�ء��\�Lf�5Em��B��+j�N9z���&=?�ֹ�L)U�9�OI�<II!_ʍJ��ORцC�I�b�^��y��=ҎmL  M<&弃�|+���%�b-QAf��D���XV��3�B-K��("g�Hm��"����:[ܫ�A����	ݚ�ʛ7r|��o��?l:2A�8���:h��{E���Rp�9������e���H��n�_X�}�ɖ�ϱp���B����Tki!�Y���Ʈ|u8"�Tt�C�z}�!�SYJ|�b�9��>�o�`;FΠ��s�b�ˇ�n�qB|��ޥ��^?�R��=��t� ���G9=	�Rj��\��՗��������B��� ��	?5��ݛ
i��nŬ�.��Z��-�#�m��r�^5��L�k�Y$)2���{І'����̺��Q\��S���e�b�gQ���CԢ�]�y?7}1�ͅ��T{`#qf�J��F|��_�:z�ͯ�)) �g�p��iH���q�9t�fےM�F�������-�Y�g����Wz�D@fth;��V����-�<�գSn&�L��Lm�����G�g��9�w�5�)�I�R��$/��kV���X���<��1��P
Q���;�:_ZY��X�ﱼ���,��H� �)W�d��B�����Љ3�ܳ�.|EZL%��q����b�OH�W���(H����`��^4��B! /5r��tw4�'+%VԱ]N Yv���)�[�b мA�a)biR�YM*�^�d�I I�M6�{[�quY�.*�-���1�J�	޶9�����G��a���3��Ϻ�<�GtW"�~��(�C�q�<s1����8�"�g�/UA4]�s�y����B�Zu4�.%<-��� ]�*����qM�w?�\�,?,��ٿ�V�2�ǋ�'�.+{��Z�,Q<�I�N��'h:��4V	6���Np--��#���;��ݽ��d�os���
���>���-�'��TN�B�_)3}u �i�ȡ�g���S�{��%�~+fĮ�+�Hm�e
��=��t���M�1a�:�G#F��ĵ�3�7{��m!+������R�ʾ����?���^_�vy
5��Y�p��q%Bq~�xW��y�w����<�F0�j�`4=��{/��wM��<օQϛ5�nı�ϓ
��Ǖ�临r��z��ĳYX>�-%���nɀ�~��T�O��od�j����Xy#����_��x�"A�?��<��k�~p97m����ґ�ߒ�Y��$�1��'���u��dX�P�A���!�8�Fl��A_��z�<��m�1�j��T��e��$ߞ�GeiL��	҃d��=��m�����J���825�1��m�/��,	]'E���*8��ս����`��Qc�/7��6������QcyiBј=��Dr�̧�Eb�Ep�c�ﴭ<p�!�d�'V�.�D�#�kS�P�%�y�a����������=9]����K�>P��:x���K��ŗ�� (h�3����*�C��T��[��Q@� �
��3I �P(߀ឨ�WC������mE�]�剡��Sp��Q;~O�1����y�-R�8Sk�eS���?�6
�W]4�Vd/,?z�Z���%z���Ttc�r9��7��x���<y�泆�I,�9�%���~ `�7E�����0�a���~�0C2��|�ڥ[Z ,������ΰ���I����������^��,�e�7zC�3����˽t�F��)5���'.��Y#�btjx�ڨ�.₌���w�˖K�+���
���=g���jN����	�>�*� ��$��Ŋ�6ҙ�ƻz�؅�B4�^<Of9髝�ޖ��]��j�e��R/\���ba�[��!U��6b�ρd_��sN��F���f'_� zrK^���_XlA�9D�Z�B�1�
�.�{P�bu*�4=3�]o�}>;��R��[����,.���c)?A1�&
I��.��������	aʩ����Ϝk��:�6� �OKvX�ՁW��R�ӻH�J�n�V�	`{��|�O"[�ݟ�T�Ť60�X�1-2���ݪ��7[km�Ci	��ҝ��.��������&uD��!Z�C���ܩ��-���rv�'��J2����U񺒒w���c>�v��*0�z:<�Y�~�	\�j��
���ch��pZ���C��A�y	��]��ʮ�Bh�6��xrg+�$ �K��t~��^3Le��m�RR��S~	�Ƅhb�w,M>rE�z��}D1cVQOŏE�$���1~�(N ��7�>_�ၨ���9��;R؟�����'�dhH�^H�^M�|�t$>���Jh�e��� 
�w�͓y�3����X;��4���{�ú����V��~�:]�rŽ�C\Fσ��DP�P���I>��[�6J,q_����G�W�Wܫ�?їm��쐤w�H˭�$f�(��-�<��`�����W1k���l3z?:���&���˥k|/
#�5��4�O;�<��7�)������c[_�pU)�Xȫ���)CB��rA
���j��m�^�"�s<:���6p��ʏk؏W�8��&�Ҋݛ�-�������Sf�FA��� ����$
5�PA�m}��ǩGa�X�E:ي�-����^�-D!��T)NT�7|�Lho0���Gv�~�=��:�0)f6$c�&���xn *�Bl�i�#�MRQH!��G�z׃�ԡ����w�.;yX��]���t,�`�1`��� 5���u.^�� ���
^�������+��:~�Y��hd���w&�y�����th���C?QKf�z �iYQ�7?����ו�o�(��欆����b��_��t��,'�cg��x0����$Z�P��������?��,QtBQKA{j�j�Q䄉d����9�2����:x��{�� ��
y�榔nj}ں�ha�̕?�k��nu���f�d�?�q�F]r_%ڀX�@�A�$n�$u�.�l�o�K���=*w�!x��Vnd�˓n^	�H�A�6u!"���LS���d�k�x��I΋�9��'T��V<Vӫ�7�pR^C�[)�v m��ԐS��C?U��̒�Ô�MY'5�Ң��Ê��L	:��D�w��O���H*- ����=�*�!'W�
@�ӹ�^�nmQ75UD\/ӊJ{VJ��;��i�Qi��m�=,I���u�����[<n<$�ț��t���KB
Nh���R���kKb߫ ��0.+4v[�%��ʅ8��OCq�P�x�t�
��M08C�#Px�߬Ġ��ydc6R��~$rg�� 1t������I��)Jq*�ǽo���b���X�9-*�]��>:��=�	yш��_���v:Q�4��S��Ə�X�6_�L_ߗ;R_1�%@EG4 ��q7�?]OA¤�ZV�;jӠgmrI��儋�fg4O��GGXٔᗬ�Q>[o�8B{~\��>@k9����V(� EcF9yp���Vз��w�3Ob���C�z�f9�����M�d�~���Ď��_�,ϲ~7��ME�xƲǘ�5����i�	�O���hO�5�}��*^~#�N�c�r�_V}3&!�<8zs�"ճ��A,�s3��}���{����:`iG_�\�t��.O��J |�qD��ۼo��<�����S�rC�N^ꐲ�5�DB������0r7ݫ%ь�!r�?��1~G"҉%ct!��~������g��x|ߎ�?�	�}����d���p'M�mg͹��:8Ȱ�[d�$�;XQ6����fL��=�iIN? _�j=�pR:6�ד�00���fQ���5w�p���h�m���|���ۧ`��8����*��Щ.�ڿX�>Ξ��t->FM��5��~�W�FJ*M�W�w!���A��B�Gqܭor�"E'�U��A��xe�)U�ȑ�Ł�m�bG�s��yvz�t3.LC K����exy��(�G�U��Ga~��#�F�Vl@�gk�{� �kƅv�VH,����4�st�nƺ�x�[�����j?/�P�{��k)ё�+Ĉ���X�pO����@��� pt��=�\���W�y_c��@0�x��e��ܺ�`��I��9�~��a��5<S�FCHy�309ľ��`��1�w�b����J�?����{�2[}�Um�w�P�#�k�0�s+kZL����rmn1 ���ÖL+��8�4}�W%��\�������KD:���Λ1Z�ٗt����߈Jz���@h��'
-�t��=b�6��5���@+I���Ch��#�}o遫�u��;���M���3�T�idi�nb@����=���fJD5�.m���*��^�e��Ж�OBI��X�J��0����^8y�_A�<�^TP@��at,�D�:���L��ԑ�ቇ|���\d�|!�u��Z�$�D6e�R�G�*HN���v.)Se R�^<0��!P孏���>��侲�%�:�P��*��P�K	E>�hі~P��4uN�Ȑ��z�J	5�w��{��;��-Hb�[WW[i�kϯQ �c��5��G���n�s������VO����;��T^ N�E�V\�(Y::�L���LJ�V)��R��F�� v�����!��͕���ȼ����Ж���m�ca������>{>1� ����YM3��=�Baj�|��0?|����1���8y ��,DF"��+�YZ{A�{��(��y�4����M�-�������:_��Ă�/J����X��Y� ���
丵/��]P8���`n88$�Hъ  ���A��7�?��F��^�l�y!�+/]��Fßu�7m�>-l^'s�ӭ�Y���~�2��ݼJt�Z\�9q�r����/���5��K�S�4����x�웎�P�)/���}'��|��`���� �B�'��Y/��	[>d�盏$�7���W�R,+�@z
8��>L�ETX�
���:h���'I��f�8�����[U_��l����$�&�_�gKr"}e0���84�in9G"o�f��7�P|�̀�`�Z{^�rئЉkT!��Ԍ������Y�';?t5˖e_��r��܀%19_�P�,�j�0l��),�_�eZ��6a]צWG������}�V��C�X��c�m$kx$�>�V��x������P��q6��z��)�\��!Aފ^�d(V�.s����L���ԢfK�jw�= }���ஶv��{Uu(�(c�������z�"���t��"X"���X�[��\2�d�uy%�);�@��UTĎ0�t����'�d���A"�]60 _9;��P��%^���`+���ݠL�Y���S���?mُL�
GW�0�gFBd]\����ԁ�v�B�����ښr�.���(�m�/�Mt*�\��k�<��nؒ������C�2����Q��y�,Y�.R�Bj��恶�|�A�N�Z6�`x���M���7�([x��>1G;Y	DF���R���[a����t����%A���֢];�B��8rGxsw�MX�^q��}ۻ�,��b�'��Va�|cFrf?�zk��H0b8��\�Ts�7��AQԜ����֑�0o���'@REL+[<[JA�D�d�<v9��c���1W�~���z���&y0��%%һ��$P���������^�m�l��`�_a�@�}���)���_��	(������|��y���q�qw�	��Pp9�F�6�Y�M�*��a�'��8�v�%�){��B�L�Գ�m8Ɏ8���
�e�0м��I#-��`�@��k�F��T�`(�WI)G���2��,��ڂN���cj_���T��4o�Q����Yj�0V����Zyn���� �4���;�¸�� ~j����cz!�.�4�4�1%�����C�L���n�&��mcO���7�sSO�v
#���ӥϻ 7S�1U=��z���{4|�"�e�C�ZgmG�e8�. �?��aF��O^�����F�cOY�CQq�6x=�w6-����O��?�Ux�k�|�VH��6��,4k��P����uv�FB�����
�ORR���(c�~�љ��P�� �'�����Ҽ��q0�&�潘��W�Vߡ���z�y3���\�*Z�7�AW!��4��η2��v\[�4�x� ��j���!�gE[�#'��&��`�f�@8��L@����џa8n�끯�{�����Ʀ-2,�k2=`��D�ցE���v���E��'8�q���*���Ť�w���
��$����R�c��WC2C���O	llҘVr����\��������=�T����].��m޽����$d�m=�6HZ���~�[�D8���a64	?�n�A����Eԣ��!&-U�0�Mu��_O�]�$�,O���fM�O�`���2i�~7��(wI�F;NЙ�7������4�U��+��\^���d;��^�N��b��v%r��Yg'(��6�R���j�d�w�В����MMh�2Pյ�R���W!�2�?�:wC+����`d��b#~�M���(t��S���hdņ�9������i�"Z]?ǰTstV�l�_;}e�a��p��Ѥ��O���A��g���xB��>fi�|���;�Y�}~���_��E��it�ϥ4�{R�����3�@U�ڄ�0�P�Ŗk�w��� <g5�s��,fSK�<)E�r}�5�,ݎ��lѭ}��*�]f-���I/��U/Ɯ�����TT�	�79���B�K�2��
�e���\���o��Z}-fǱ�E\�������K���.�۹�)��(�Z���@�͑i~�i0z��(M��C�a�<�n����!@m&u#}�1��z	1��w�z�z]�2#M��j�g�]�B+�����;���")�n���?�6�ȷi!)=v�u@��Ɗ�۠׿6 �{V���dB�@(�e�����,�g�/$�,�MN�0|���!7۳ӟI�RR7��6hK�#�t��UvIlW<)�nZ|z|\��-�eL�t��_7xaEj"FvY	��[�����;���b�����!���+F�+I(�N�oDc0��,�^l�@*��G�ȧ�\������6 �w�H�ǲ�|��)ZQ��Q�|�B�k��we�����O"r�� �,���p�k����eA�स|~����4G_�{���Ж�����>z~)f��l	K#�9�q�)��OI�*�+%ψU��_��A�s��L'�V�����
,�u�2��� +G�:�ɷ)~`�SyRZ"�}#+V�����<|jc*q�Da��ڡ�����w3�]���ҧ��:�B+�x�w�����?kn�
��6���+�*�D��Z��@���)D����8N�c��L�1a�8�'l����:�|������*�m�De��ͭ�Ϻ�I��6G+tv,�[����@rW��:ȷ���,�������$���BfD9��L�m�"������(~��W�y�"�\oC?�U��U3{�����$C_R��CD+Ƃ��3W\��\�P��T �X�}'�;�	��V�x�-��c��9L(��ZzF���y�����t���x7��C�d0񱊮
B��-v�zkg�կn�*a~����)�ƶ�Sl|{
h�ϢDq�)7�υgY�$2\����g��x����Nu��-Z�=|���zf��d/>>�r�4=� ��p�6�}-��h���<�H�z�tDn,'���:�8:�ͻ��3�U�M����
?�Z�3�^�ҦRR�+t�ϟ{�^��G~�:q��b�hX�`���ˊܜ���Y�b���,M�|y�����c�Q�4Jԃ��@�њ���,��u9�*_�;�]6ޣ|2�"m�
�2�7�p��j�w�>˲O�%���(ګ����}�p�x��� EON˷����y�o~.�?�TebD&S�OE�<�|y�_�e�Y(E`��/T�@ow<�ϯ�tPS��#��� �\3T�T����J�'$�3���X?�^#�hAB�d�6��b�p��7S��AP�7f�9�\�-�8�q���u����jQX���_��`!q����O��#�>2C-&G��Oa�gF⢠B��#[�.7�����l�P������ �����G��$IIb�U��}���b?�ã���Vj��j�g9Ch�ΏO^qa꿅�M��U�r��F;�,W?t�9��q�E���^��KM+�C4��I��x���]�>�åء�GJp.C�M�F��țZb�d0���$�4�/���U��HB7[��&�~J%ޚ��2�8!t]R��܉R�����?�a�!�J�s��ߧ;7���5\}��X'?
���ƒ��`�p�y`Q4��F�.E�i�����7(�B�jRfK�A�b���&V7���o�wQ\�ќ��t�1v ����i2�;Ѿ��/?�z�1��Y<��'�e�t����u\
��I��uqN��x���n#����ז�!�X���� ���ql��L7j�\/u�~��<��mǯ�@t��3�3�>nLF90������a��+'r/2�m4�[!�r1��U�At
B^|�D���TNߨ���٪�@��S��;z����Ü�O�RG��	K?�1�rjR?Z�KV%�-!�<��8"���Yvl�k��
2���HN#�?)�T���4�=�r7�H�J?y�E��<�M�3��S������_�.�9)��L��U|G0\&�8��n�m�O���6���W��b�絸9Z[��V&
���܉O��<n����i�X�h%��1К�LOh&k�U���c�`�;$4��'PEz~�<�8������8?�Wa��{�	$P�bG4܇�"��Z��a�� ����.z��EC�Q�ԫ����._�i��Vw#{_&���M��[�qȜT�M*^�:Ӯ�g�7c��8au��(���ּ��1��}t?C�j����7�Ak_H��h#c��U�?v�����c$�Cם�Zht��F�U��`#�'k{������Dx�8-"���|�YN�C%����a�eo���`Z��[/���"�Zu��N��]6�z5�
f3�	F^>G��O����Et�HH>�ۗ���]�H�XB�V�#����g�8X�]�L��%�����(B$�R�k��:�5Oz�iռ|kl6L����QZ۞�RѪ4��Ѱ�j*XlxVHYEB    76e3    15a05| YI�5j�지�ͩ��9�@P"������KBV
-�@��)�YA�[ߒ7ƐV�>�f[+X�*�G�6(3Z�bO;r|O�Yu!��>,4�N�CO�u�;=�U���h��D$E�W���H1�4x|� $�+WQ��Y�Z���w�������w�ԌxZ*�R4���.b�g�c~T}я�
=��>�)�փBb+�����O�
����|k��iw�$Ai�'�X��b�na��h5eƓ7�@gS{ؒ��c��1��3=���u#�'�����l�ȹ
h��葘�k�����''�g��Լ[�tǘ�|�����Z'J�Mc�ߞ�4���� Y .a��~�yBR����2EK�a0kb�T�!�d|�.��oݘKc���ٟ���L�ֱ}|��J���8�K�Q`wS�m�݃!P
G+�CZ�Z�cꀤ�!Dհi,3����Y͗�\ӟN�Ӊh�������/C8�<t+O( YӉ�f�Y��`�!f:���(��D!��8T(�@�Yb��)T��KΨ���.�{z[��|��l"z��tд$>��R��L�-���;>J�G�x�eK��(��ͰCþ!N�ߚ�46���T�-hj��=)���u&}iF)8x"A������ĵ�|)M2�Z��-�{|��ٽe�+_�C�?K��[>M�����dҺ��g%�;]�6�i��hz����d��0��N�kc�����+�1伋7�Re�ּ��K�4�'w���Ⱥ\�p�׀��n��������4n��+&h�H�`��N�F͋B#�'B8>�'%ڤ�(N�� �矽�c;`�x���{�R��Ű#�y9�j���'h5��8q�A�зHD��G#�͘��N�A��v�Z`�e�~j���ZDyʀ�
Zw$����_t�b��|�)�R��X�Dy�f���p�>,;�[����5c+ Q�0�\^Մ��w!�2QD�$������SC��Z�A��/�_[\�ʞ��(�nb��]ʼ�s:�v��=G���>t�΅�0�ݲ�����W�>yd���b����4�$C
�f�ǊQ��v~2W�ǚ�҄�Ŵ��B.D�R��o�~��r�Z*DTF��0p�GdB��-H������NҀ�[?S�+���J���K��˨�Et$V���g�Eqc-�j���3�_�[{�Z�7�lK��7�Q��o�� �*v��'GU���Y����@��7������f�N�
�QrPO_E��)m�,����@��1�7�]d�~�h��� ��R�ݎϮ�Ѭ����V���X�����_>�-*����P�Ow�.I#]N�$�݂��,_���pN��Af͜s:r��-�|"�1!t��{ �W1��\ǋ�LK�xl�菑�F��7�T�1�W_�
��Z���!a#0/��'�Ǽ1kM�E?�`S5_�5���D�{�?.&S
I�Jq�B'�.�2��V�z�Ѹ��T�qe���"_�>@��0LD�����G�|����/��K �|B�~4)2@1G�v�m�u��x,XW�9��4�u��X�a����m�l��qBDnG�kW���J�R�zZ�~[T�3�K�P����T����A�-+c�´�T�,�D����i6���D:.��`�g�	��Ѓ(��[�k�`$�\;�� ]"`w�/�w1��v䃇y���OF-1���M���)��yxK&���i���?�.�)8�����@u�l�-�1m���|��O�^������F_z)����m^�BF��v���l�˥�s�i��q��+�Z�
ٯ+��u���,�.gk�B�G��25��4�ԔWL.{幱���m�����;6լ�p�^�w���d�IB_8�C��g�U,ѭ���Qޘj@d{��\��O-7��b�z�g�r����U�F>�_�w��A�M
�3����
�N�,���F؜O����"\��0��J���,qрd�	��q6l���M�.o�>�� �������+>��s���KN�˧��h��3��9�@#�(B/�9�iɞ�E ���� D F����\�Op<	�@��k�M���&9�{���D�r��u2gY�bVLh���%C�r�B�v@
Vz�Ud�}�TS��?�d<���΂�	�L�綁\����F���W$�Eq��Ƞ�B������%ؾ�%v�	��J��+�JV�-Q��qh���_|nGA2��1}t]k�[��&��K;l0�C4G� ����u��3[�/�	�F6�<%$:=۩g<���ϐ�� ����@M҉��۠�ژ��d���M�x�,�@�΁f�\6�[�@me����S\&?[:^��?Y�ڙu8cn��@?T�@t�/���q��8��R���A��I?�f�&�ti�z+���< .��\�����B��o��"��)k��J��˨�m���[����W��m��<�D�`�~��d����FX�]P)6�#]��hF��^�ٹ�,АAC	!֓Z�F�OR����=���'oέ�!���w�Tc!gZ�{���B_Z1�m�jbP���WA��� ۪���麼�xu5_��
�����?2���>���	~�X(CBOr���ݬ9�ʶ���]��#}��3*�r����[� �f���`�V�?�Г@�ĺ�{��FL~�5��*=���C���6?�H�Q.;��l}2�l���-H�_}|��/�Զ?6�!�������",���)]��x�W\Wp���f�&|�߫�:ܬ��n>	8��15�(�M�Bh�����X����j��
Q�V��w��vP�\�~�e*A�pLOY�h��V5�2�J�~�_����'c��B�U�DU HSS�>�U��1>-�TO�O��9|H
��EiKj�H��t`F{-��Pd��q��ZT_�H����Mf�ck�h��jrR*K����z��gZİ�|YEn�6��|G�=�Z�0ղ����[K۪�/V*�����ֲ,q�hd�O�i�"A���A9#(Z�r���
_��	&y��ƃ���w?��J
q�|��&Թ*]��� ��q�9�"���j�*��L�3�&/��ۨ���$�J�o��1����F�!/�w3��-}������k)��qPٰ�MY2dYΠ��!f�/n>{��t�/^]�1~��;���-@��CU"4�-|�U�Z��SLE�JTn�����`��0`9A��������	�)D�޾�?��o��B�}<6�5|�G�w��+4i%'�{N1��$a.O�Ɏ�Ȱ�N9��H/䲁�����v�6�h*��H��j�Y3̰�{T�B�4[9���8�
g�a�`��/^���	?� %}�����`��R�of��fEt�����c).k*�`fY���h��;arnfnJ4���x�meL��n��4�dC���.u�Y�x�e��\�1�SML�~���������𔯞����ů�4�0ʯ��t<yδ[-��@J���V�f/�2�H84ˢG���|�w�X��y1���F�����,���^D�NN�둝�ܛԌW��M϶8�B�ʾ�(��?���_)hL��t%0����R�!��/�������c�U��I���n��1O���9Ma��KF�vK	Z�("��X�͇
�a����|[������6'<W�50�*0�^�h�O�򠙹l]U�X���<���@�{,b[���ǉ�kd\İ�	ɀFh��;�΋'��p.V�5�-hps}�1�80 )TW��y� ѪEl�P�����;[&HU��@4{+�j��:�t�ߜ$�IJ�V�$O8���4�{����т��S˄�����|%�{�U)/Z�m�e����v���D�'*{�8@�V2j�;�fwI�Է���/���0�d���)���L;Y�3A������=E�z��/�$�l,����n�]�{��C�d ��S5hn<i�����Ή��� �__��s70�jͬoDG>��Ts+�p�NΰQ��8r�Ir�{r�"L��!�j�]�'��OG <�Y���&�!��00Z���
��`����J�p#�qSh�@1WQ�Ky����}#Q\�Xlz'$���uQ�+�*5�zqϴ}�7w�S��`��y|�Dy|����<u\A�?�B|!}��ҿP��$�.k�MR).�Wƌ?�d�l�D�{�u�M1#��{Oqk��J�(�,�"]T�5t<������e����,�N�r~�j�Ư���O��FOj��1�Cޕ�����ݧ ���$�X�<�S��	��&O{R/��qWe/:c�3ss�g���ʍY[(�+=�N�.,)I��<������2��4��r�1�a����m�;�k[Q���	��7ƨy�{y�\����Y�5"�Hӫ�F��VxU����%�p�:�gɗ�v;*g}�qbj>'�ޚ�8>���ꋂS��~��Q�V�6�����g�(�[O�[ą�C�'`H�_��C�����fχ[{��3�N�T����������T��mz���`��I��2�_�أ�7�
dg?Qh���&����`��Y�
��C��l'�����wj��e���ب�Tw�;`�@Ӿ=�Ww;��y�Z��U/?��{���Tie&���z��i���N7���4�䫰�8�s����jl����b�wv�3�y�jcPJ����q�,8�ME	iU����5������P��G��CF�:�M���g�#KD�1����W�C����2ݝE?��S�L-֯��8�.�#�ۻ���B�$!�h��m�SkS-�^��RrL~�:�H�~;�P����Fҩ��c/������u�!W@����Hu�ж�� �� �.�%ނ��(9�8"��@�(��V�V�Ii��<`�{�6��������F'���[xC�� S�C�=���H�8�)�3���-�u-M�)Z�4	Di,�S�=�+���#^|�h������g�!N^���R5�E����$�z��ueF�`���m�=$5}��M���G��B|~�7y��T��d&QG�ҕOK��������,��H�����>��_�)��\&%��%���/K"Ӿ���8�
$��	얥X���'
}/,�0*�W���'�����F2�ʮ5|E������ű�391
7��b��M����C�|kp�!i�
�ŉ����+H(1aS*#U A����Or�q�:����C���o�� ����)�G�Vc:�.���Iv�j����1.����Ec~����-7��"2��Nt�%� x��[��@&;t��������C6���G��d��M��Us���~��
��3E�ݕL�q��"�s ^)�N���v��sI�t���E<�n��K2��jk�~O���p��795���_e>�u��7I����x�u*Jb�+�ۈv��`��\M�˦��Y@��ZD1�T��6��ƭ�D�Ɏ�UG��oCG�3