XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m}��B��"6��K`���^-�6�'Q��]d��X�A.����[��i�=��B����.�(�V:���<u��qϵ�+�#�y��n�I70��tz��b����l��E�'�f��%�&�=tJ? �hך�������y�Q���;f����߄�"��_�^2�v����k�&��X����!�3H�	O0ȩ���/dӕ��c>��?�6�{�������^[ުr����s����J���^~@T��Mn��<4_ɀS����ue� R���%�c|�?���-C���T���6��o��w+X����&ytzD����?v��ߖT���W��,=Ӊ:����#i��j-t��w�p��ͥ�Ǭ{@�R���aH�<j���.��>D�	z(�6���X�[lX:�PW˄�쾰1M���^k��~
%1pXU��,�:���R�����s�wf��/�c���_�A�A+�y��V)�g�UA*��D���L��a����m忊rkQǴ�ƶwRx�$alώ�V|G�$ǣT杔�/G�<�>$��Zʩ[�סVȶ�PF�-=Q�A�Ek�=���C=��>Y��iBN׀��$��5s���:/�7Rc��"�@���.!��stTD���؆���?� ���ʱ�r����FK`Q��)}�D��q'�S!�9��7Z�����=?&Vi��i �l5r�]	�M� �3�`�5���|c�`�0� �|"XR��@�ڎQ[�cɰ��};�Y4����XlxVHYEB    248e     9f0�'G�� "�<p��	. �8�����J��T�o�����~4_!��ASBX��s���� �R�g�|}wt8DO����.�7��C�6���A'Yl��s��A�O�m�"$��e$��!��O��eX�ee�������8�1��}�#G�I~B��"�X�i�����6dB�S~[����!��K'��;��LW�۲\�ٴ\�9z�l���%&J�+)`�*�ሳ�ɶ+�̓zL��+����	P_�`���Y���嫍�s�ܧxs]�[�b�^��U��m����L���3��=i� EO�ݺ*gT~(�9��\#��8}�3�����B}�Ҕ�~��U5��-�+�UҮ�ۻ�褋�?4!�m�$���%�E�
q���;�Q���ʵ�Ź�?�++n0/�Hf��[�+X`M���Āk����w,A���ܢՉ�oTb �o,��4�][,�[��s�8��U��)�=�|�r5ʔf��9Q͞���,�ީ5��"�e p3���`����QL��e ����>ގ����K�s{Mcs��	y�tDW��6C9���\�WZ��k^#��r8��-��.�����5��-{��V�Pe�v��1�M�_���Ͱj_!��3G��/Q� 4�Ӏ1�%�Y��i��k���/���β	=�{2FYxW;�:��{+�O��ạ�sw~!�+7;z ��Sq�Z*I}����Psl�,$���,��"X����{y؃>��g88��Pjt��y��X$�P��#I���P����� ��)��۰l�m��]�ŬLTn*�~�l��喥��|=��b�$����--U�Ⱦ�3.�J��lڗ:d�)����cF����$<�u��>4�o{������I���N~1)�"V�с�5�&���x�̈́��j)��X�Gp}'�=q��	���h�U�0H�0��	߿��=��u��쬡�li:94v�0S���I�O�����f5�P�.�7Ŭ#ڗ*��}��uAz������� �ؘ�k�q3�4Y�S�Y>�+X3�z	HO�*�-�I��O�D�S�&ޝ�1�l��D���2ė`o<]��5ŔA��~΋P��] �aM!M8f��U�r) m !��������ì�!��L1�fi<�+\����~���?aC9����ƈ����������1�W�K��D�tŀ}%�+�[�,K���A�%"̄8U����3���Ͱ��e���M=���T�5�ȭ��3�ßȀx<Z
p��}�,�_>����#�OI��d�H��{X|yE��� q1`��S��0�(ճ{�n��-�BN4	]F����H�<D��*��	L��� K}<^����j�o���Ū+��>�PJ=Ȍ̖d��9_�?P��Z͕21Z�v�v��0��t������g�M�����-	#�VtV�ؑ�N�N���Վ�J��;o���Y�y�z�j?K���������͉sKl���i�Q�(V3�=q4�88Y"�͵��~z��z���z�f�q.�����ѫT��iE&���&�>,�;��JOŧ��(��zK�(���� ,�B��//Q"��puW�B�M����E휠E
��L%�mNl���x'�
fԨ�
�?�b�so����cnY��9KVs8�����F�}�������H1��&�̀.�N6�ݔٟӜ94�ӰX�t}�Hpw�t�\be�f�Kq�A���<g}|�F��m��:�6�Bky$T��'�7�+��h�w�P��/����*���֔a)�WdZU��1�_��gtG71�]�
I���ђ�7`_��j��zȣF��%W�v��-ٸvõl�M�z������H2Yۗ=���[�R\j���4x�\�V��o4!U�[�=;�i��W��|���&��(P�t6�ǔ���" �Fe"�@�\��F�����*/!9sjqe��fy���B��t���[u��>��%Q�5B=�Di��38�,���7"X��7m�)��=Ks�*:�< -�q%�E�7tՇ[�5}S�z��T�lL�xGD�X;���.g��];󽫋_��hB�,��u�"��Ɇp%79et88_�)���|����ֽ��hޞo���|�Ҩn���q��N�K�r^�W����@|׹�V��7�m��Ə9^ Ė�'ߔexD�T�#�˜������5���@M̞��H�����u�(0�G%�N�v��)�Ȱ�q?N'�m=ĩܝB�>���2�4=�y��\�� �ؠ$*xH�W �I�S{�~��K�wT1D/��H��I�q�߯{3�(f��kO��Ps����b�h��m��4�%!��b��-N�N3I+���̚~���A�B&��3«?��p&���h�`���*�h�4�K�͍�Wa<z���ʾ6"M[�kJv]yl�<]�r�s}�,=�ג���}��^�:��FU�Iz��`�*-���i�d8e��ѨJmO˵-�!N�+