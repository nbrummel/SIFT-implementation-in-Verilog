XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���?��n8�ˤ	a�ф䊯��ӒO�\@�aF/�Ө�?�u�_�v�˔��4B�'� ��`I�-c?�D[�}X��Q��B����!�\~��&-uWlE�	"�GA���G$�]��-%ő��kV��J2V�4�GG
���Car(�]�ٲ�x��9��.��Q�$��_���IX|Rz8�5Q曛�C]_o`׫x��5���	Έ�@H	�G�~�z�]���n���I�g6&�[m+� ���y ���Ol��9�a7�E�")��P��|�`�����$Ԡp�0:�*۪��${��i-�"�TҨ���ܿ89����y\G&�)�5��n�k�WH�M|fK�V��7�g���tq�Ѹ��z����I̧�
̮�W��$X��5Ϸ��m�db��P�\���/9��D��v�>��wD��/�@̝�4ABZW����C R'��!���iQ�d��)�y�=�Q>Z��������ǥ��U�u��2��Z����Y#K�[-v����6��͜��������C��3��#��S������1�t����ʅ�zxp�����'���#A{�d�v7j�x�7��%d���_Ƞ�Mc�{�&H���q�N�b�Aޓ�$�8�D	��;�ʨyl��G�@E\d&t��͔2�\\W1�x��_-�yT2w����[8��K؎r��>B����o�����b=䣗hZ��O'ٵ־�LCy��T�Ղ��u��;�`M�9���g����T�!��?��K���I�n�f��բXlxVHYEB    9193    1ed0�qǴN5�*�ޤPɬF$1�;��m�Z����I葞s0��1�j)|�H��YܤÌT��&=1y�>T%T��K� �U�%'-�.���R����Vl��*�� ��
1��Z��x�S/���T��T�'��8�V���Ϸ�͸��p$PO�:�,�q§a�"�\�nZ��G8�)�74[��e� 'o�V�U=�w&G�D\^�V�5C�a]����%��caJ���a�d�.�\R����E_��E#)R`���W�A�':%�3Zf��@�~Ӏ
���'�'�U�/�6��K<z��Q��q�'qu�Q�A%.�2��Z� ���wH"|K�T�Gȩ)Y}ܫ��HQ�ȸ�.�!ӈ�F��ŘL�i�<��L�ŏ5����|��<*�h��<��\��"�-j7����e�H?AF���X�]�)]��Jv{��ᣫ
�|����B��n�%��D*ʏ�
y���U�0
Uuo��_���`��r�S�@�T;������'�	�0�#��!�s�+v�&gRP�H�砧K K�t�T9��F���8��s�Bt[��_UѨ>��<[�YY[F�=�CC?#WT{�ZX��ĖzÙk��t�I!;�dA,��"q �P�i��/�L����Us���tmP��$��U�2U+p�/rO�h���z�!�?��R�G�Rl����}
�D��~g%mL��I&���H/kY_X�!ѥ4~����Z���KuY�sg�Bh[d��W������A�)CBI+����̺}�w
���Y����^& .J�ݮb9J�I����0 _
=���Ϧg�n-�f
hi�.O�P	3�������kcW��1Q�d�a82��E��\F�����Kr7*=�x{���~;X�#*A�Ѱ��?�3��~=���������g�v�s)�{���aW��ڹ��+fS�O����5/O J-0u�Ʀݤ?��9�'��@J�(��J�.�1�i=�%���}�[�L<ul��I������j#�Ӱ�I������j�~�g.�s=�\�O�[�!^�zQ|.�I������Ǵ�oGI�K��`���p&8�8ݽ-h2�-J�G��L�_��۞"���E���G5�h�!�������fe��E�iMNl��[�ٙQ:��Y�=rT=����ێ���*{�R4q�w?;�;?>w�hҰ�Z�|vOޥ���%�ЎaE��"�5 ��uh��K�險Ӝ�˃I�ݞ:�:�@m��l�
v�-p,��QyU\�6/!�|T��%�]�K`wMJn�jP�0���Xܝ���cc/O�J�A�\�+�a����%CL�:�!8��zQP��F�f�w4��λo"�s�F�ִ��~��+��`�'� 	���y#�Q��!R�Y�N�i X��� �*�o��h4-S�X�5c<C�8�,�&1�Zg-����;�k�Z�gY�3Lu ��j�q%��=����)2.��+"O7�O
T�!�4?�g��$f��?���u�Ō:�3�)���$��� [���}�%��s|�6僊"r���ͷl��Z括��_3����!��<���c2���"S�e�&��Pn0��+�Yf�*;��*!��{ɞ��������2�,�����b�0�`�N����x��W�9����H?+��,"���;Eh�����g��ފp�W9�ÙN��to���(�2(B�d݊��F��w�w}�k�FW���>mw@p�N�#���
�����N:C欮d���B-:|�BĜ@�;ܪ�(��~*�`�h��d�r��T�\�m��9�߽��M!53��d�¡�<��H��z��	1 ��b��X��mw���`ٵ�}ۗ��y�V�c�ۄ`\Y_�JC�f��Z_C_D����o��H*z+������<By�H�X�;0���*�1��W�B�t���,�5��Ő�"����.IB�`t?ϝs���}�ͩ���	�a���
��S����WZ89N]GL�It�}>�w:���oc5x ���"��v�F�H��#r^-��B��[6�i�z/3�=�oan3ygW��U�J��2�8?
y@y܅��,�B�U���_��R�yA���F�b`n�U�Fp��Lɝy4g�T����/��`"��:�!�R�������^OYB���=�)W|�͟�I��T��-�j�8	3
�`�|>�B��űaW	u�*�ˉ����%��4hf~��LW���5�;âJ'���2�P!���� 8s:��A�U���n7�K�=�P}�8�"���,a!�|�:�%�m��$%ٕ�*�)%T��4��g�Dc#�-���k����S\��t���|��+�œvH��:�	�w|�d�h��� .�뇫y6��T��h�,�J���a��:6�� �:	g�G�[`gQ�2.�H�W^�%�k#ܖ�Cb��֠�&����:fK,l�f���@��l�N�%�f��93�S����P����7�Y�h�̟�����'e���4�klA�E���6�6���2�쪄��Ь�L^�Br� ����ӿ�%P�!�9s�t�p+t�T��. G�D'�P��֨��Uf'Ma&����v4t�oF��p��m�@�+�e��M�a�뇽�ׯ��
;�B$wZh�k�ϟ�H]���~��%~�L�;�]uc�o��	��y�ӏ�j�g�����ݵ���(f��`z;���쇿M���䅶�J��'W���yjjD�*ٸ���W��t������������|�>6j����k�Œ�%
���Ԇ'>P4@��~�l+�(�̄���5a9JL�Oy� �I��/
p����=6 rͣ[%�g�B�J�G�p�6��	Q�p���o5aGR���S_	h��������S��V���;�����R�2����j��n���0#+=�/�}�������%��*}���|u0�5].��&nv�7��g��̆wsC���K�lȄ 'iTsw/W@7�︦}��H�ؗ4��݊��Q���*������>�W_�bMv��E�p�u�GQQ�1֪�&�9�Ȅ�pY�EԢ/nSjN�C�璑x��X�s0L��	];\���o0�i?AT/�奜�VW�c����.+�0�R�*@橺ݴ�_g�Q#��V+���Q�O����1�^/^��0�מJ��W��
����!E,`9���Ǧvؒ������/��P߱n�1�������)����R�TN�N��_|kX�;^�AH���~wA@����Ľ1i|��4�����2�Y���y/�A��K��A �� h@���1�G5���_�3���, X���24��u��֮󧼪��}x�>���I;�t�.@�M=l��p�)���� �¹YK��Kk��Y�3�K��4�W/g�?WT{�O"�|���p_+��.Ǒ'��H�v�ۏ��9��S�1���Bz�v��u"��9��%��Qfs�^�@L���[x7x��}�h'�p�{��1�>�eJ�@ʗw�<�[5���u����~,!%u������,���5���T���C �F�P\� xo2+��=�f,I!P�)�%���-�a*���j��Q]\;Wrt��=ZB�U�
3S�<�$�[�C�>0%�X��.B�� 6m�~�N�2דd���*���[���� �-�~�u%�w��Zh)s8)�I��ٽ;���'��ўk0���I�k�0�hn��"U!W�|�U���+eS�Υ#��ܘ7��I�^ݬ��gt1PW&N��hK����{�ճs���	g����
f��I������?mK���ػ��(,A�_}T	�,`�1.���&�n�ɾ�~�#���k0qO��9�P���	�>�NRc!k�8�-u���� O$�aym6:�k���̐��b���w��6�X�F; ���5=�#�P������{�V�ЉT�GWdM~��g��Bl�	a���V�yPR�B9>v�&�����F�E��->\�G�n��A�sG�1.���|5�xQG&1��+"�A�u��%��Âtk/���9�gb<��~��@����M���!�*�堒Rn��j�9�ǉ��:�d)��My0��tT��ů�^"�ƃ�r7f���j�a��ڍbu �iϸ����֞�+�/L�������a�������)��!v'IH�g7j<	nFi5����c���JL|GZt_��� �s�;�*h��͆u΁��,���*զlܻ�5�p�������u�~�-\���q�X��A0L��W�Ga�KM��t��F	s����g��5�&s������O��H�3�"��%I� �π�)S�������x�:=zl�&���J8G��6!�e�����5��Cne=G̸��$�~r��Q?0Qf��\ڣ�h=w��?��q�=�78H3P�G��ѿ��@xk!f��SW55�~y�"Q;��1?�y'�,~����V�0 �);�^lN���Ylݓ�f�8c'��M�ƒW����S~�8���6͓��dp�ś9x���� ���A}5�bd,(3�Ǐ'K4�!y�7E�E�<��w]�Z��������6���]��XU���X�Iз;�]S8I'���,�,2�\�
֐5�=��N��)��xS����� ��1���Ê�J��BAM�D!!9aK\���%��g�Y�?u-ԲZ��Z�L��@	YQ͌�YBC`k�OPzQ ������{�K����aTw���f�>�O��u#7�{��+7�����WNc�����A�6�]H�Q]%�ԫz�cҔ��>���l�yh7\K���>`n��t�ڢ�'��`��L��/.;{.T�� qӛj�Z��������gd��d�ZeY�)+�����L�)��#�~�(+(���Wbb�W�S�+�X���+�t�K��Q<�XWj���Ir�
���=:��֧��˘_�� ����(��P��NB�]��B�#��<��̞ڼ�~��oZǐ0��O�e:��s��Sf���j��Y�G~���;�H�UB�2r����a��ܤ��I�3^@-���c�ݏ�x�#���������?���2���m�Q��D���p�z�1'a./�vڶ��9�o�������Sf���6�֯<J1pNc���m)NѪI�(�"��g~眑m5FB39��z,a�7��lx5g<�K�K�@�]�E7��s����.��Ac0�Qꯃ�ġ��D�ۍa�?���?�	6k9�鮃O�FN��Y��	>Mk�f��͙∧��/��/���B���ò�B8 zA�����$�q��nV�x�@˗&w�b�l�4�XE��=�UUGf��k9�B���.��l�ҙj<J��w-/;Fw7�A�����GQk	�Np�J�����t���,0/_$���YYȋrO!S2&�%��t�ZZ?��?�V��1�[�'��U\���J��(�D���=d����Us��M�!���Bn]�n(���8C��c?�ڰvfF f��[N��]�勏z��$�#׮�t�bkO���aa�'��	ʝ�S������/":@rtɣC�)0��ݴ�ݝD�'.2=�PV��S��_5�^�7��ԙ6s�W��V����sF���jwW����%+`�Oи<�q�ԙ�E���ͼغ��e��<L[��A;�f��&���R��&�0�ZVׯoD�}f&��c'��Z'��(RIx$���U�=����;�J�Mތ��87�q�|�ΞR0Af�[��~�k��2�@ �Lb<��K&50����E��)h�ft\��%��5��<޵��6��>��`E�)A���J�R=7x%_���`�r��tF��
б|T�Y���SR��쨋'Zkh�M���&X��ѝ�؇^�b�W�-a��d���71�Q_���V�wl�H�]�5Z��h��0L�/Km���d����,f���X*i��@
��AJ6?�u3L���~�'	�OX��l@�}AxM��JV�I��'Z��y�fˆ��a�������i�L#���O�i��9��M��Z&+�N�P�xoxY.�jB����Q��.�ڻ_��g͓W���-�����Ե�d#z��ꦍ�������������O���\5��O]����b?�1:�Y�3�I1N��a=<+�Fho*�E>�Y�͕�}o�(���ƭ�oX`bH)ğ�/O�/�U�y��_�����Q���q"����k���EBυl>9(t�.]��y
#�
�%%�R�K�LD_A6,�w��G�"���*���P;�����>l��Pt��w��������L�>��Sc����*,�:EF�=�Vs<M�[,�E*Yh�0�}��yzo��&gͣ����4��se���
��O�)gw�#uD�g� -&����V�Ϲo��Ȝ��v��i���gl%b�$���3�Bۢ������wG�G���`5^�PM��\"	��V!�Xܻn&,�s�Ǘ_&h9HXS�Ԁ_]�i����9�}n{�KR(O: �]��[1x��C�x�s.S�N'���C*O���B��~�'*�F n�������A��tOb�Ej��~�XTM�C���)��|ƃ W�K�2�c'3O��$�۽">��� b��xsjj?H�ʩ�,rP Y5h(κ���F�V��gk��%I;������_��@;�E��T�؜r[N��-������ r�&��K/p?.?�ϣ"G"S�Ae@֟��V��֦\έLM#��U�mh�;�@ ��?��q��n��y'�(1��jZ�3W�=m� P|�>/Χ�dP�=*_V�K�v|���f�x� !N:�	��	/G+�����p����h�ɩ=[Z�.8�����97x�fdez?>/W��_s��(>F����/}� ����[
��K���s濇��:��_����B��b0���a	ҙ@��Ү�R슌/��-;��3�I�x��>�Ϭ~�^���ۮ�9��GZ��ʔEz��.�L�~ع[R��.M��m�������(pK��,E[��09�7�#�n���	�w*��=��7*(]�T������Zg7�C�5�8-h��AJ��`|���df�1�F�pJ?j�T��j���`��?--:q�X�._�{:;��,�U�T�����mn��==.�-nA���T��ˑ��ex�b�pY��&S�x�tc��$�!�p9�/���`��T�ks�
�e��;���R�^�&%˅����'BPL+���� �����nzL\w�x�&�)��j��0m+I�l�ݥFjp@6^�K�,T�50�jُM�}ũ��b>����a(�7����������M�wuTNIV��,�����V�߽E6Ⱦ�4�$Q/�v��!��lu���б	�|s���o��Q������r�L1<qK��';i;	���v�ٲ]�,�[7#J6��I�k嚤R�|.s$��z���nG�Θ<�P+�
�s��J�*��*0�� D�T�!�e���`_�Wc$��V8V�+~rF��@c�G�u���,��=a�N� ����ӿ=q�rw�\i�%#��n�\����C
8΋^�w�Y�N�Э�Y�i����|U���-���������;��.��C�Z �ksX���r��˴��1�<
]���	���d�di;���t�]��s:]�QN�o)��%��9�5;�lw��P?���N�-.�|��[o�m��uG�`�D.؍a