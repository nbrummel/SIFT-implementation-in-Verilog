XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k�H9/����I��%D���+b�$#���PP�S���Dn���S�uB��Րu�N��Hzr\�?ɋT��v������2���a5#�$MF3�<(����?� ��;�Jpۻ��%��?�!
�
��Z7:�/dˌN�S�j�9��M{MMj>�"W��Gb`N��� �?�� 5�Ǿ��ʙ_M�8Х���/�æ��m���!�@~�YoF=�ڽ���>i���Dp���U��m��'N�U��kb~���y��6XC,-�
��3OX�����d;`[g�A�e��Ew�Eu`F
2A<�4��j�B��K$���:�O?�CŐ%:V�Xd�D����� ěvd�٦9����~q�3�=I�E� �m���^8��[k��o�ހ+�P[��2�}�K�W�]ү�^��kϼ�����DF2h�`H�6h��3��SE�Kb�4��M�gi4���Nţ�O�	��B?�=���1X�M�pzXyb�����Z��Ԭ����f���)���n�^4�����6����Sz����U��%��|8�Iݒ�o�S��gE��iG#��=�?�J����OQ���T�_���SN�G�\�L�HuҺ�1M6s;0I�U���%��D��	�v�W�\ï�`/|��L�"bL�ڍ9׈��8�lLjM;S"Ka$rL�I�2�(�/;��9�<s޻�:a��7������܈L�-(��=),�\eg4di۟��rת�˹ק��UT߁Ll��cevb�VXlxVHYEB    50f8    10100�ds�@Aj�ev���>�g{�hC<����,���sk�)x��4��xk���m)H9��܇�ل���R�����eJ>AS�����S4̜�A�E��Ҫ1)zK� `	B₝��Y��4�]}�]�A׊��"odl�P�ڄX���'J-��>H�s �T���lH~�>�U#X�9D`1L����!�#H�A���laE���V���Uxb��'���c�L���X
��R���ލ!M����Z�9���f2v�a��t�Z�\S���Kʁl����-�]ڽ�a��ص��E�oLN���	���Lv�LH��&7��`*�R��S�Ϻg������F���R�`�ުދ�;RJ ga^�,.ah>�-���&�hY{9w�K����	���4?ʴ4��\'�i �$�����DH���Q�j(z+@hl�SU�N&���Vֆ��ǟ^��,��� L<5�"�u�*�m0n`��0�u��v9�m�W�B�?����.��93�~//�����]�Z���r���N�m�;���Dn�M�k��;N�J�cK�ک�SsFzlF3 �G����I6��hJ�.�
L>����g��o��QR;:&`P���8�����3�^Vj�ZX�%Hʰi�^��SL���<?�~�Z:CV��Ox�:�2YM�z7-�T�q�|�V���,�T����SZx��� ���.9ЌU�2n����ұ���kK�u��[��GJf	Q�M��O@lݖxm���k��ܸɎ4��l���m�	��]@�WL�@cS+��;��z����DP^���� �"T�j�ڠ+*�Be�zX
ₐ?+�����t,�8u����y��S�ênc��5�
8��������x�w�	ܨ�e�(܍Q��gA��dh[��G��'��N7vn{2r]�Ʉ�E���'�>ve�:=��A�?iʾ��F��]~z�Va�
m<��z��s &ѭ�6	R��;!��xM����x��o-�.��5
O{�d�F�=���:��A�b������%	>t�,�`J�nfL�[��� �hﱥ����f	2�B^E?:�������8�"��/�&�=��EY�B%l�¸��s��e)��]���{�8NV��Y���N2/������>�sz���a�$uTG?9
!x�Tr�k�gN�ݨ ���N�D��_���;��V���A���y�Д茊>n� 'Ȕ\|�UWV���m����B2�x�N"�n�bԬA_�\��˾�����Xkߌ����Y~���3�t����'�o�ep�~,uU.�&��T�R��ʱΏ������o��dA�Ck��.�`*�ח�;��|d]z�P��6�����ܷd�K�{6�τcy�51���!
�ƞw�o՜��~7�H`��Á�U[1����ǄM��v [K��<���ክ�H�ӛ��YtBP��Hfp�f�ܐ{d}Z �X�dӛ��
��.0�%B���X�`=w�����	{�~lm��BJ_���?��cV�ݘ��I�)]"�Ь�/���Q�Riu�<�I������J�]o%]
�La��nR �HKz����o�O�k��-�j��l����q�3�et����e�[������w���Aj�g�s���Ɠ+�fY!C��ݔ)�`}ͱ�AK0x^�T�
_�܅F<��YP� ���:,��N��q
kh�$���v��`�E_3ąfqiZB�
��SS;j��5���w�&��Tĕ��x� �e^���n�X�k����gᎎ|J=�i�q(�$[q�ۑ#&�'��ڔI����df�^�NO�J��T��9�+���C�֮�"�O	½��f&F]���U�@> g\�U��60D����P������� +p/�IDC}p�Gu��O���e[ �	ʵiw�����]�~˗��8(�H_�T��R#Q9�����d��y2T)$�x����.�?�p�*V�٥�v��.�~���J����&�,�S�ܸ��Cu-����R�[����B�	&�̾-��ʵFE!�%鍻�h[����V91�b�G"�ȳ�'k�ZU��.��+t6&�8Gz����v�ZFz�%l�"�:(���NQ�{VJ�h�V��C#Q���"��	'�����+a��\7��tU�����`��}s�a�9R����Nd�������H�&��5*�b#Ľ���$�j�J�r����#b ��F'l����l��X��s/H�Λ ���Z!�o�.���;`e�%Tݔx�{2È�Ol}�?ĆR�+c��2����%�\d��M�&]�a��i�=�!����oM�<�\�o�(C�ѫ͉�ڲ&^+�,�������;`��G*|��tU+��R�-����������9��l���v�}�$��hэ8O�2�a�_�Qf,��c*^1{_����W�OX��ٓ��=��K�ť]�Ԯq�����4݊�oDO��=V������̈gm���t��^�U��*����?�/�����e��K���g��6�LY� s�$e��j��!�u�%^Zo3�~N�Wk��]��H|�������S�.��3K�6��E�\\
��"��N���8��~�!<�ܳ *{���5&��% �ՠ�i����7
x<x��AoN X��_7i����rpJn��$�il���4�]��O��)��r���]��)EJ����[�j���H=�k�0g&�K^�(5�u�-����q�!�"'�75��uSb�T�Y�^��U N�`��9�zkIi��pw�C���tZT���t�Ћl�:������1�PI:����P�u��
�/5S���/Άn%l���7p��2
D�������2'���-|ݰT��D%Z��b��8+�1���v�I���=U���2|֌������L��`cf�S8b �`;�ϒ$)2��1סLׁ֮.]1��tܧ���w�����u�T��ɑ�u˶��I4�Eŷ�J]���@��+,'�f������Xv�ԯ�9��(H
���s涽�Lw�a�P�w�W.�g��G
�w.g��L���4�"i�~"o�E8���*q�]���w�=ϭ�N�/�yD����y6�V��7IPV2l&ٳo��G/^U:3�T���n��g.GN�@ۗ� �
>���	�[C��$�ܑ�HH^�`S+@�~�z�C�w�\aQ�6�	�q�\d���(�&�������Kv��#%t��h�/��m˿���mM�@,��8��� 8a��qߛ��2���犢�	���<�d'QH9�eh5��g �����B<`l���7+ӷmr�ԙ�0�������Sr����G��.K�� -G�n��܈�{��#�L�0zќ�9@,� �J�����
IK�>�-�����^&e��z�D���8�DB�Īq{v�-�ߘ�έ�pa���]�i����:�R�}�!�K�ꖎ�q^�:�O�Xj��\O~�S�!�<]Ld�;i'A]��u�;DU�r(�����k�I�j�*dC�RN�w���s��Tw�	�m#c�d�d��?����!��7�xDR?|&�p�:���[iQVǥ���%*��6W�F���\��%��p�G����xŋ�B<K9Y�Z���o���H{�)��1w�y8�ӿl��]r�XX\֤�e� E1p�T���*�~�
a���-Y�ys�T*ܟִ6D6`�5G't:6Đ�����t��2�����\�����\��M��ױn�+/W��!@�)(Ȁ�8��T}N�&�9׫�LyN�B�+�:��<m_闅Ƭ�#Z�M��o�(���4����-,\��8%��x�g����Z�� ��d0[�&Wʙ��Ѩ.R��o�I��R��BO��ʼ��i����"h[T��\^�|��z�-�-�^�h��"S�dD;)("
�e%�6��$A#�L{sX%
������<`=�Աꭓ�Y������
V���p��>��;H��	Z�u�,������W��hL^��.��