XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6���	�������i[�L��WG�"8=�0�-���o�6̠5Y��;�m`o�nL
�s�����YE�&O�v�_�?�6��ay��a�7t�cR����#�"3��n�TAХ�h�`i�K�7�-�0c�O������^�P�垭ƶ{砜�l�;�����v'���W �G� s+�`o�'���Wl+���c\h,	F��ϬD���+</}��x��T�z�s��A��zup�~$�F�;C��=�^�GW����q^�LE(��	������J�2R��UI�	t�RG)�g9M��}�X W�",
��js�I�Krp�����=BXe|�L���a)Bࢮ"��$�>�y��RʷIޠJ��娺ь����"����sd4������ܔ��F��(_V��{�7S�F ��*���Ya��PSg[����ct�V�m_��^�W��t�:6Ԩ���t��ń��c��ٍ��',ɮ��!t��NB�Cg�.����t[��J5LE6��`��#�U���e��r���e�H�KY�9������W��O^��L�ڶb�J����d߾W�w���ˑ�k��b��.{v�y��u
�J�e����u=9�$�a�g�r\km}��q��e����t[�Vߙ٧��0JY 
4��P�5�I҅�&P ��(J���OtQQO5�*h4�s������9#��.t��2�t5��$�j�1�L���[���p��a����`��$w�9��62�C�^���dטގ��Za5��
o�XlxVHYEB    507a     f30>��6kREk�Hڜ�`��d��SM1��b@���k�@ÀoAIʪ�����7 ��b�5�@o�wC5�i��м�e-�lk�s��U�y���$ 7��yҭ�:T!����R���!p*(�J%���Lrw�[�� Td2�A%�Ni��0�������RE=�ό��{5獤d[�ޮ2e�^�+]aWZ~Q5�%�ͱ�3XW���K7זw�K��=3���+)����X ��߄8�M!���1�[��<t_�4��g:��'��?<t���ϛϚ!y�-�0@�R��ʓR���Y7�	���F�A����hW9�5yFG��A }�,I�|�E=�1��?�Hs͑v{F���V�E���a4y��X�W����q��xG��.iaB�J�'!���x~�����Hx���N�Yu�Kw�Ls�֍	��.o���,}��\���mJ���v�;S���lIr�Z��8O:��������']tٷ�&��/4k�]�&WO1RJ�1�3���G���;���HF�.|F |�sW姷�������n|Nr�{��ҧ�����.I)����أ 5������L��h�Wk1	�V�I��N�l�;(�h(Z�t��#�� ��2yd�%C3H�vh�>�qeM�	��j�����wŃ�+������g)�YL�,O��v��^*��6����>�M6��e�S�8�ȥ_�-.�Q/�&��I��GNs���|����pY��fZ+↡{1����̂\6s`��B'�����.`�'��S��os* U��T��+ M�/�B�St�S��pi���Kh�c�i�h�?J���3�74��tK�Z����#%����/�@`�� jw�1�/����!fBUHkrl��L��8z8�v�J�w��>*��t-����I��DcP3>-S�Ϣ��ф2���>B��&��O��$�e*C�!��,O=l�%�)��AX?0'��a�?yVA�)m^��`�E��s�B]�֌��R��n8ް@{v�Եg���5�}\dM�M�,�rρS��q�%����Q� ��t�w��JP]�i�PfgQ�Z�B����kK��xQU'_Z��0R�@ �\b�Ig��F�"G���Ԙi�v��
.���v��X�����4�R��zȸ�n�ܒr,+�F�-v��Cz���ډ�H_�ή�uȐU��5p�f�G${���z)p_)7�ka�1�)������?U�P�߅���cRӬˇ�C�ҘU��������={k�<�wlyۄ�����$�&DQ�޵j�9Ap�ld���ƻ ���1�������m�8����B��>���h���>{��v���/}�#Όs���}vcso!M��A&5�	R첗,\hV
���Z�S�)؟*�8�o�	U�DK9�ك�7p>����H�q��$_�|��	���;#�����5tB�BH5#.���R��L�D��l&����oc�ǳmH�� �c��4E��Z�Yk(\ku�
�]ן/��õ��I;/�w��]�ր@��Ď�c�1�a�]8�d6����1��VN��qp����GT�$I'�`���7wh�<Z3*��.f�G�G��K��hw��Ǖ����Q�B��ЀA�|�I��$Β=W&�X����Iy��]<:�G���eXkaVCbJd��9�R�z�gZro:��R����L��� <���{�(�L'��=p>�J,o�̇E VOLsr�`���#�'�����pKy���ԹA�G[*��.���jBǏ�5�ڼ'e�ʒ�ԍ�r�W�p�"���h�]�B��R��8�6�"�_��j�{e�c8�Cv�t,	�aV"l���>%H8S�5O��2t=������zmQ�E�բ�(uK�|������ZT�ϛ���s T���{����d֓��Qчߕ|�n�����?� ��eeL��=ma�2�6�D7I6�<����O�9��uW�/:D��ڣwV�w����6�*�R����Չ�+������!�\�����������:j���SJ��4ʋ0���,��ALb�����L�]s�E��%/�[gW�L'õ�_�8l�����=b5�"c�\čϕ��[��z��.|��-&#�w�у�n��33
PN�?@�
���&���?y�?9�9���Pv{ؚM=Q���p���ށ���Gb�Z�;S���8_���@ub���!{�����8[ݔv� 0�V�	 Q�`��A}ĪzR��Q{�W�x�,� ��'�H���5،��s�%{�VB�c>�lF\;�ta.��C�m��Q��]�q��� ���Q�E�`��k�7X��,k��ŀ����`p�����r*9�!�q#yRX���B 6�e2�7$��*tH��/�N�,Re^-�?�cc�hl�Ĩ9�m�ؾ���I��9.���x�Ȫ�D�#o!���m���� �N��3D8ISQ �O=�2���Nn��y�CUd�e.���yj���ot�'W�-�?(���';����}��f���!�e�Y>"���~�[M��e^��nf�vka��$�������v.㠗�qפ�R�𰻇%�wq���A�K�UK.N����	�0�=Y���Y!��v�Z�	�g�۹���b3x���aM>#�T�cZ��w�)����������ɔJ���<#�]����U�&�
f�9�SP�ͨަOF�#�r�od�/Z�k��vr:b��!�.l>o�Tԭ��6wά爟Z��.}����g:͂��*<�7���9�	Â� P�s7#1�B���+S�;���kׯ���C�E���h3�q󝭆��5��ȫq�Ka�!*����8=��)����OV(Uf��l��]��i�{Х�0"��۰�]���Ҵ�Nt��B�t��5;4>㒉%�ch(���^�q����/
���L��{7j��BM�$'h<fΔ(D�I��P�N�?�4�q/8w�����
���-��t:�%W���:�Պ�*1�a!���}��~�)k��4J/�����O$<u�Xp�� �2O�Y�)��m��şs���� �!U?եu����"��A�n���ͼ����=v�_{��wD����9��v �'[�2[3����'����텑���݀� ߅6y���_��Bi�*4��Gkw��9��:��&#9g���m{�%{��=�pK#&�æ吿c	M�0�����^m��b_�"�d�{^�Nw-�{/�����J��Bq��銣鋣45��e�"M|���>*t��=>�i���aG�U�R����TH�H�j�q�������Y��"�+�+?��)��5��Xxۥ�6�6�o����Q�:���b�-���f�����p�6˙�,�q�=;V\�3zQW��U��p� �<��)j�LX��E���pk4*P����=�,�Y{d��̃��n��&�l8�]�&�����>P4�#ྚ ��r�TP&��'�#0�E�^��H	.��3o(��;;���������9fӆ���x&~�e�*��B�,v��V<vH��a��5l���J�'��5��7�36.!Nv�ېm�v���=���Q?C�Iq����@��no&?�=��ɰ�xA��31�L�}Ur�q��`����uؔU"r�����2:~���i'�bԖYY,���v�(��$�f��"\Wa��%D���zWrY���L���Q�Q�U&�l?�b�L����
�����!�-��5��d������IN�!�b���!�N��z�~��<(ǢRشfO�1���LT^�r	��X��u�f|���s�?�ry�2�]-���p