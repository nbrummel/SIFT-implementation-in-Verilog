XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Y�s��.��~] ުjṈ�:��l�Rf��~��h�yv��')?�)g�I�"2^����ZQ}Ϗ�DBX�Ǉ�R.���c���f����HL�t�Lt�~����Pn�T�ᛯ���k�$`���t�(>oTȆ4*��Dv�{�~XK��:e ��7�h\A���� B��Hk
q�F���n�,�5?2)����P)_U��-ET>���B��c�m^V� J��z�=��9E��:-����Q�u?$|ud����m,��Ҳ�z����'ӳ���=>փ�k4%�U�W�?Ң�:-�ќ�*��`\Q���tR�ɝ�����֨R�w#]�V�=/M�@m����6�MO�ʼ�X<�ao�+/M Sx���'�)� ~%g����h���6����a�S����� ��,�����m3 , ��f{đ���  0w�o����ϣ��1���vhr5ێ-JN�S�8���;���+f�ve@�Ā�Ze�g��]8����4�8�7�X�32�|W����qW-� ʸ����m�Oi��
��Q�+X)e�C^��D?�U�JD;������dg��0�\���	���(&�om����>�S�����b$�S�I�Tb��9$VvCX,����d�0i5kX�*���,&�iM�o�����XΏF $15��r�c�jN^4i��-�{�p-#�qH�~��q$QG0���
ǜӄ�_(Ң^�g���O��>�5��?�o�n`ۼ����:�9@����_X�XlxVHYEB    4a7d    1090��Ej���-�[�h��'��C��^�Ě�`�nv6��V⿵��~�"g�wn]h�NR�K�tY0^���# �te ���ΤC�{^�V	��~c�b��~�q�vn�Y0,��-���G>��X(��PO'�G`"�"�?F��/.�����vI�����l}�!�t_����7�w�$}���"�9�" ���k �8�N�d��J6tpT��ujm���sn`CF0,�aZ.�ɽ���gz� ��8��Q���ۇ�y�����S��zQ��e ���&�H.Ʃ�A�rsi�cQ�_�A_k� U���(ח�m�Pɿ	u�hM�L�EGH�@O3��5�կv<�L�P{�Vt���A#.ueC��*ϻ�~]Qp���2�h�9�9aܡ�y#!�	�.[IQ��iL�'p���Oɦz�����+Ca<�Z���Pa��հ����w4�����vҽ��5;�$Qߖ� �)���{�e���V�w���]�������@���>[��4�/���$��a	$7��
�`�GD�x�)����$${Yᘇ����v�pe@s�x���݃vM���\��A��ל�%/�GM��,F���$����)z���R��E�Ӣ���2	�������Sw��90ܚҢٹ���2LQ����{����7�@��']>�a���sX?-�6�zYk�)	�zJ�S����%�K���Co�_�]�9x���$c3��DS��!��&v�4��D�4~�.��VH�ŋ^�,���W	Q3	�%��a�3��B��R�wX)A�Q�[��3�ʎ��|>E]_����3}yoPc�9���&��C^�۔���ӡ�S*s:�M*�`Di��4��Ys/��?�)
��4}������w.�m|����V�[�%����2"^
���6��`���������e��U�㡐�iY���ə���<����"N�z�a���t���g�� W��\����E��8{P�ccY��|����1�!�=o?�2���������X�ڧ��,�v�Vމ�J�<�U� Ç	��9ٍ���J��}�z� Z�����|���N"�A��n�B�����߁�B�N-�q�o[�W��Ťл�T�b�U��Lp�M����c���{y�xq����^w��J� L��[���n����/@��.�M_�TXQ��w�����6�2��y�Ɂ�2Y�)��d=�­BtS���^�8��b��RL=�8������E���k�d�Zt�oʫ���W
x魅�e.�adxުV��{�Q=�Gl��kW���qf��p���IH~�)�_����2�>���vB"�n����x+��=�SB�:$������OB����ai���B?L��W"�}�T ]��p����DD����yh�!Pj��TC|S�l������:�����z�0������u�q8���U��&^�ܥqH��O޺�1W���iI�A�#�z��;hq}/2�Ծ��cxc>#����h�w�`}w�]Gr���J2��D�[֬�?���2nS
��{�"O�\��t�0��y�<,]�aG��g7�L�ǣW��=V�!n)�\Q�Օ�����gᎂn��d�'űH�w*�<h���
��A0F�
���6S׾�Ǔ���b].$ɹL��K�����h3l�}�`���Y��L������{e4��<�J7mRp�(Q���u�(4y~�iq�a[@j�]�
G=��-kz���S|��Uw w��	�F�WĬ\��=p�J�[u��R!˵�;��g�O�+J�ĥ�I���;�W7�C�MThL�M������d�7���j��� Ǘ�i��N�ƁV��ѡ��r�<�q���:J��+����?S����۬����v{q�r:��9YĽ���H�ga�F�0�`��-C��2����YB�L��.� �TsB�wgz������(&�������gj�z��Z F+�Z�i����Wޯ�kX��Q?oS��mȅ��p��C�Cԃ�b�zO�D��H���~�A��~V��m�m�V(��
,Q�D�*t�a�E~;��x��{��=#K�2J<.�Nt�C��#�c�M9X�`��A��^4�n��b����t��Hv�/3"'nS���p��2R����|{�2�儺c������S��<���R�4����)�����{J~X#�����ﭢ�Ǔ�@�ۜ�V�H�H
��*�):͌z䕃Jៜ�?2�,���x&�'R�~h����F���@��a����]R]��3�q�������c@&Ltd���D��Sl�'�3��yF����o��LY�-&r]ɪCyݳ)Y��-�V=�.��Gܺ�q��bw1F� �D�>�0�/�%�����`Ulz�0�D�p�2E�d,�,�F)�ŏ����]�^y�"���>H��� �2T7���@� &�����h���3�$���P{���W��G��@Ų�lF�ѧ?K�g���m�fӺ|�#�R�V���,��vC� ��z�3ׇ+;�Y3w�C[���ʥ���B��I�����y��C�̈�3-F7�U��%@�wu��Vh�r�c5�avؑ�|���T��_�+8M�-Cr�Ӆ�J��'	��d���p��0,�TI;��^|Nu.Thyy���1v��&�L?2t�=�GN�2�������3}'
*���_1v'�huW>��w������m~��9��sؒ���1�R�@�U0��B"�NU\C��-�% A�x<�*f���������O�Zi?�'j�f�"1۔�w�Z9H�?����F�Z�"��ڠc���T�G#'��#�D�
NB�8��T�l����}��Ӂ�Q�:ⵓ������3�&���6a�5̬��'�sj^�Kw'ѧ�%�M�Kys�D쑧%ަ}���	��<�W&k��RC���DO�zW���9��#���$b��f�jT�#:��^nl���B5Tb���O(M��J���ɥ��	N�z	#�_:����I�/׽N�,�����l>��9Ș�����~>���G��^���b�Vb�v����mMd��<���9��{F�#����WN�xC3����>,��Є�2\ɰ�/��r�u�e�������p³�!3�0���h/*׀�>N�#}��GɁp_��@ҽ�R))C�ץ�v�G�Fa�L��I��a<p��#]bK����0� 	����f�j�Tʫ�\XVn	�Z`��wA�ă�*<�V���1M�^�� A�ar���T��o�?��NG35����X���l��=�U���A}%�ńH���^�i*�w�)����g%y�9^.N��zx�_#�77�4��L������%�޷O�Hɰ?��m�x�ELg�1�Q�4��F:Iω�����q�#ߠ$�݅W�}�-η��{؉JU���$1��(�0gMu5>sv��/z�5욌�3�V�.�6��l[�\�{�$"��օ��=$�8��:f���҈�����ۅ�w�"[����Lrۗ�W�U���5����b�%S��j9;�&.y+�*���)	�����H�x����ԙd� 0+X;.��l��?������P�W��L�-T�!	�`�1����w���Qn��V�ؽ
K��G0a�4��>�nBYh���v5+���m����#ȣnmw[xKYǷ���$��L���N���������ٖ�Ǫ��Q�%E�~ *�HJ��'�Es|w-m=�猺��릥�j���	)�0���
��y9`��(�S�_4��J
k�2a$0O9�a��y�h�|���'\%��䜲�-��ۜKD���:k�7�2#��$�����WA�TT���1�0xXiG_NJ|��%T�J�:���P9['01�Hu4ů��[�qz��؁��8
��K�휹��O��b��Ef�0_$�xN�졔>b��P}���w��W�Û���Hg�p��ƍv�����%]��7�e��5��u�yHE��vK��+?6ondy ���=p,b7�c,�tՠ2�R�#���h�ӷw��y.|�چ�(�%�HQ{��ot�g
M  �4.�j2�L�V�4b�l�EW���t�}�s�Y�ȳ�^���S�*l�h�!���M*3