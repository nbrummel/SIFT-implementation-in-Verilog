XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���T|��[�C��jx�,a�&�4u�F��n­��q�a�x�j�煻�2�����g-��[�EM�i��5z���OaKԕ����k]�R��"Y{!���	��a���2��W޲��3�	30�0���,����q
5["��S�1"u�� ��m�k=�:�/�����v�9���FD��!q��o���"����z7�c;���L����n����V�C1��c�3�ƶ����Ԅ(S芝��v�?�|�;��6~���^�&�~�)�14<�q_��
��L�D�5�	�R���F�Xކ%��y=�)Fn=F��=�i���zq�NS��*�=����6]A#�뗼= k&{Q,�=y^}Sըm z{��cd�X���%��{���9'������֌G�D���J��=5�ǔ����=���Rm
��u�k7"fj_b��M�7�σq+J1�w�N�CD�8�}��Yh��nNሻ��%liοd����.�-]v��Ǟ@
!a�G}�gO���w� ��UK��SjH:'��>t�OjS\Ő���r��~nU�o�:�K�*CT�n�o�s-h ���1Ik�X�\�S�U�V�2����:�W���5��F�<��G��gr�x��
���bpf�G�4`��g�CF/�d��رC���ǃ���\i�
M5Ր��a ��}p7i���J�|����b��yN��@��' ��AR�|b(�s�Y��"��`���p*������Wa��F>3��,#z�)=#�M���8�XlxVHYEB    ea93    1880����#	��H��4�Iڡ�˽ш ��ә�!�"+��HuH+=Bc�B�X~�HL��Cg6�\<�Y�ė��f>���4�e��^.�Ҽ�^z��<,���F�	�3>i�;�d����e����
�6{�;�S�
~L�*5߃�E�I��&1�7���h��7U�l�Q�m�2����
�t�qA��M�G;zBb7�B�b����J\�JM�8ɝ	X��"*���0{"�l��g���q$n�?\l�O@�#'qvXԍ���ɼw F�d�?D��L)6�o	X~1/��?���B~����{x�˰�4tE+�Uf�� v'"���nV����0�4�S�n`[�ӳڬa~WQ�r�(c�d���m1z����$�7��}���i���B�O5й.n}���Q��nl�u|	�8؞�U��;4��袳
�g�z�����J�f��ȣ ���D�,cȻh� @�.H�����.js�T�PdP5A�}�#^�4p�(S��ǻ�h.梹�a���Z����#�=b���������Ϙ�z۷*3�Q�5�?�CکQ`�(^�׭rD0g�Qnl����w����������3VE�����:ی�ƙ��O�G	��l���"/j�s�u�|��"U�⧲"_��:��0s�f��WÎk���Ǔ+�!�/dV����R����i���*?)�7���d(�*^�Ɇ�k!-A��|��4E�/w]��w�$C(��\'Pݽ������i�@�M���:`��鳩m�+(����t*K�0���ݽT�d �r� $㠔�D�(Нe��Rך!�[��6�J9?��Ʀ� �>ѳ�F�&tq1V]��OX�T��7o,�9����"s���ߒ�W֚��Ō�����q���)%G96G�"�OT.W������v�e�D�/C�$��r�7LbQ	i���K����A]�a�Y���.��`lL�X�ٍ~9�Kͱ��t��3k��ãx�~@�2x����׮BǞ���� �g�e�#�F���!�}0�
nW�����'��U���Kl&*��>.�>�qn	�4�L�?5�
�+�nM±�'��R��7�!³�zV ��WE�����s����ͯ�φӉ��u���IeQ�?��5�*��幣�G��l���J<b�ck��0U����2h�
9�jO�C]�5��,��_���4�Wdz�*%X�Mbѯ�����g������N8X�,w����v;L�B�fPQ�rq��j�I<bsr�NͣW�0�\Z���w�iE���+�q�ޚ
$�WU(O���lQ`!�����|we�g���6��{c��I�8B&�\`f��L�Q���4���d]�}�"ӊ7-�'s���c�V J�qWS����4|��o��%[e��$�Hu�r��S���Qc^��˄uZg�s%�O�6ۃ���:��\�����*ðg��3��n0�Ë_U~���rx6��q׷�΄� ,'�Nr?L>��`⏂�. ��Z���ӿ�*�^|v�����N2����
��Oe��i������H�%�'��?F��|�7�-k��{�PT?���Mq�c���ni;�凗˟@�}X_��M���8��4�?��q���^�L�	�Uf[����7�M�-_�m2=�(�l�p��Nf�����V����}������c�P�V}�F??N"�bV����d��� �v�u�e�O��!����Y�pA���Z�PUP��۩�UQn-�f}������r��I�A�2���L�:�4/��=o�V����4$V?m
G�hv�f���u�@:�yo�1`���k�|�v�=�9g���M�����c�B���u�h27�7���+���(T�	��	�V�"����QM<����VL/�����p���`�X�^ 6�/�TOo4n���o*Ou������O��Z��C�[�?혽5]�ϣK��*�O3����l���H�\��*v�9g����'C9���85t�$����>i� >P��ڔ>YMv�g'�r��A,�[]IH��9���^��.>�$N�������� ���Z܀ѩ-��>���k�h�E�5�����(~�-I�+5�#l�#K���>�(}�I���k�n����C��E�&b/�s�����eП~ߵ�8��80,lx��
%,$�6C��p����E����Q	���S�*#�Vd�.�Q�#1�(%tI;W @�j�����;���K�͕7b�B��_ɟF����H`͛ª��I��*0�V䤓�ҡμ�ۘ�����,H�;'�w�@���4�aAU�;������P���K�*UB�(v�wf�9A���4&S���vr�SL�%C�\��ݫ�����C/�n�s�y4�&(�Ż�� H!o!�_:�d<�8a�h��^;�@̎���:&�C�D'c[I�p�^~^y{)P/�ʮE��$H���=��6A}�@/RA����I����>v%�C,�H��tm���{x���o�jXV㪈4�c��>�V�B���T68��:���!�ݤ�忐�&�?ŕ�p�Oʈk�KG菈�'�Q�*!�"e>n�֟)��ss��б�����շt!-I9��e�ν �6l�Ì=�e����K�������ǝ,��d��I����XAK�ɴ�9��t����
��~�g�Vw�~�5뾙��M�'���s֫�	N��B�6�����^#���2P�p>e���VȀ�pB��dø5�&��?���^�8W���=l��e�^/e���4���f7�l\�t?���qrY�:bT �6�P�W��d}�Op��!/*C������~b1nW���{�	2Kw�|B*Wh��˨�TzV ���Ւ�x�Z�_U����j���m���Nm�"|�0f�I��.-�'.3����o�5Uv��E �'�7�+ Y@��ӂ��!��1�7�Z��K��.ӵ	Faʾ�u��0�/U�sf�(/Y���
f���b���S����ii�"`�;��q����ߐVn�1i�yT��)怯�c�g�f
�V.=���l��1�i������i��P�&Xoc[� �r>�n ��'�z�l伻�ݔӍ��]2&	L�g�j��)�h�t8@~kbo�PBI�o��I8� O�#���E\Z6,�������Z�аB��Pp��-�x� a"�h̊~�����(M��"�ٰ�Jќ�e�u��3���m�^�Zu�SW&�!��J��9a8��f��ƪkp'NԚ@1��=��A\R��V�zh�i�Q��'� G�N2mq�~����*{p&_�3l x���d�W��[55�䞫h�Y9��E��Q��`��f��e����=jI��%cG8�>;c����d�;�C�b����-�����Ѫk�wm�,bp��|~s�\=(���G`�p7nO��|������X'
�=�LY����!��{�A�'�����`���'|T]ZN�^�)�x�����x?l�'4�Ţ&A��n��bK��O�W^���2�YV�/�Tu�"n�\Ky���՘*�;?nq�E�g�&[K)�.�����A�E��i�L
�����c���y�,�`����������[���%�)Ûa�e�#���-�x�R�n�v�Z���x�3�:VtH9��X�;�p��m@�L6�GN�G����[ɥ{�0q�����7����d�8K�F* ��hB���YF0�8���[�����hvx�?�ܳL�g��f�c}Z�z��?7E�aE3xlsI-m��t/T$i�J9��U0p�S�T�{�
N$�3N�:�Cʔ�ޓ��\���]��s�6�a�Bs���VX����9�`��֞�G�n�W֒���c2�JS�.��g_��H*�*Z��Z G�������@�G�Dę��B�PG�)>�z��t�+hz� ���)���y�5:S�,�
>�`/�~�uB�7��V]n�6:��3!n��EK�Y��E��u���d鱼����}&y�R��5�%^��b�ꁇ��Z�9�9�����фdRm(�in�A��^V,��P�t�Up�%[�*'��bV��ͤDs��g�DI��*MW(;'���Rs��*ч�xrb���z(�\���Al�����A��a)c.���&�g#�V�T/.���о<�UBI�qr#�~VH�0^��b%��K���礨"�35W��R��0&�͒�c��ځ��@ "P�&�g��5������q�D�op�O���Y"5��Yi��䍞 .�&�6F�B�ze�JβS����Ei'�����̚�S��O��)F��hnS���Xj��H����J���]�=��J����1[;�W0�%��R����󿎣�H��)1h�;���Ik�y�)g��eR
��;��������F��
=��� ��|��{YH�=Hzozd��I�����J��o��˺�=�1c���[]��p�6h��w��:JH����az�2ܓయ�ɧ̿ht0V ��nTۀ6X��������\XI��º�j�6�\���>����vO�&�w�,m��$G�������A�ُ��ao(����i�Bdc��j�,�#
Ns�����&��vSi��鱪�] ��4t=�'�۷#�װ>1���8EM���e-�T$�n�Y���c�ub���
\@W�YW��t��2+���D���hAB�_4V��N\x�#�K��s#��H�g٢�Wp��h�|C���3�%I��k�H��;Z�����q�Sf�`�ɦP��NW�k@v?��L��
 �	gH��Ft�]C�8��/�i��:�;���ω34���p>��!��;"����V���쵔߉�8���ҹ)=�׏8<�d?+����J�]�t�;�?V�$�c�A箬EJ0���^G0֒�w���Jx��1���H���
K��q�;s[R��ᵯ���N�B$����'i8����.v+����ǖ�0������[欯��IFBA�@�5_�b���XD �J�z�}�������ny�_�N�����M�����o�2�K=���X��#���)x�8�$	�S�ʝ��G"�a2xC�����Ekk�6���!&�Fz�+����b��Z�.z���v������ɇ8}�S^��p�lq_�č��0�v"�w!{:��͊�,g�E���FsIJ^�
h
[�`$��E��H7��7�`��Ø�z\b���V�0�B����s��_�S��I$�S8�ݮ�ys	RmĲ� &�섞�'�Ĩ�����|(�6Z]�S��U�*���yÔ�(�x����0�E�螩[���3�U=.w�� >	Ϭ�t��qsq6���d�'xߋ���_�A)����Np���ծ⫷A� �֛�Ws�F6WN����b�j�����[��B{7�?e��;�P(������L;���Dt�_;umԺ����+�~ˠ�Ҷ�NC��B4J����M,;'ϣa�ԉE��s4,�ȷ�7� ���Y���[�|��=��O��Q�Kw��]�u7��[�&	��qqX�^�&W��r���+Wt��.KY�xc׸�J�ٶ����&�~r��Y+pqV5>J��8X�'�6��˗q慿_�����r*Zq��f��[��GSX<F����~4b��0s��NhX�V������=l�H `i�R�s�h�'q�� �L�$�����)y������s�D��$��4(�3AF���OV�cث)8wލ��F�x� 5����J��H�"Ă������|-:WV9!�T�]��3���(���������ޘ�Ö�$�y�;����T��g_�֥���MνS��
�{��h3����qWK�E�D���_e��nv��E7a�Ei�&eo*[[m���{k�0t����6��ӢSe�� ��Y��p��kԉ8�I������#�я�Ib[T{���b���+�E�o���Z3��gL��#��7�H%��JU���MN��1)x�W�~,�PDU���/�U��6̉;Yl��D���II
خ���*T���EO!����v"���t���T@?�]D�^��,�/���n��ΓJ5��=S�&:Rk����^e&�*Y��.@�zUtv�*#[w�