XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����*�Q�&�Y��U�Ԕt}��u�PAX���2ٳ�_e)W5�ˊ�~�9����`�����B\��V��q9�B��<ag�Zv�^<wFb6E�b�>��%��!����l�!Wu�K�y򁗗*r�^���C���ka��7�W��Q?g��ɵ�i�� ��T�~�-���YH��@�@�z�W�\�3�]Z9t[Z�7YVR>��A��=�#"nr'�Ԝ��n�b(�7�$?�jVڂ��bM�<(_�u��e1��}�1����vѨ�]�4�����}mfA�yX4F�*1��x�+uw��$c�w�~s��R�n9$�U�	o?b���"[(}�ڷ\�e�U��u� �[N��:p5SH���g{j7$�i���@B%�Xh��7����j[��Œ�7�$#��R6���|�a�5�ꋃ �+x�{�#�g�?y�#�Թ�z�m��y.�}l�شkE1ݷ��ꉁ��>x�����MW���a��������� �c M��`�`�6�/�	HKۀ)��:$��@G�c;Xe+wV'
;���c� n��5��'���ӹ����S������bޭ�(�Ψ�"d/X���b�g6p}��?@�sRr�3��x�K���&~���=�]!c$h��T�$����?�<�zv�]�@r@5Kx,���S4!�Cb*��$4��`��F������d(&&�G�v�15izWt@ݽb��R$,���H�i���1����E�cҙ�=��O�iQW�҈eXlxVHYEB    9de1    1670�
�>#�M��k�l�&���蜴a7����!���,�E6�:�fL��q��o���{m*�7g�l��I�D�I�@��~���������+��9����Y�Y�U{_�Gl���b��U��5��PK�e�,ᷗR÷��S��IJ;!��d��\�k��#x�-ʕ�]��Wh.tK��sޡ���i������LXw��"����:�poHt��<aA����Ln'�޹���R0
�٪� �X��#�3hB��n�~OV�"�/�_��La�~v�o��@�]_�_K|m���χ�2����{9C'��m�흛�B�?i{�c�mIf��Pc���+Y�e���`�҇�j���$��7�&6��P�ҕ<�W/�α ��"�B)������Y� �~��t�6���(��M��PΡ�˂O�����Tb�/�����<�ȝ%2�Yq����$P.�<K-�h0��s�)��Rߟ�ĜI�O�VO��l6b q�ZW�Fo#�ߖ,����s���W#����W�>;�4�8�5����k�o��� �����Y'g}��;�Z�x���l�x��ԅ�Ѧ**?���*�iNW"��~��,�->R�Z���A
��G�$̑S�!:Ӛ:O��[�>�rŝ�	*J
��X� jC����	d��~��z �L�4�]I��Y�����W�isC`~����.�^w�0]'®�U�_Av�5���A��`$H G{���e�H\ܸ�C9|���2��a�!�ϖc�hG�Xi]K�*���<�R���w� �}g��Q�{ɼ�-��E����9V�a��+����&�}�]0���m�p��s<��6m����D�>�o��D�џ�B
���DG~<��B���7'+��W'�Iq�v�j
σ`Dw#��K�̝�Ҵ.N�+5�滯��o�d�|�s@�4>�$��|��a��$���C���8�	k6�^I3��	 ۅCek@�͆��M)1ecWC���Qr���D'����D���m�)�)�L��	- ��S�LE�u�aF��n(��9a\�m1Z_هf�jA��	���[�����x��
���=�0��v�+W��M�A��$�U�+<��z��v���[�V�꺒�q�|';x��3�9�����ڜ��Jd��	f�Ώ�&�cvY��?�z��P�`��?�����������E�w|�|��e�a|6�O������n;�|&p#!콩�VU>��0{���?����׻��$��c��0V�|$�j�M��
���:������f�_�J��	��0���װ,`�D\�Q|���ۿ}Y��B��%�&i�+S~�f��m������������Z�&zC�7�L:�1��<R�^�Ĭ�N���z����С�[Ǒӎ�\j>�u:��J�x��	4�_I���c�PKq@��ȵj�}x��?�Sy/�ɉ�cIk�%&����LXmL�oU�:}��a�����7gi(c�q�5'�v�c��6+Ofn�YL�cE�v�9��IJ25z���]B�3ޑ��i�C�{�#�c������Ƶ���2�I�N�c�FGt43�E��=
^�S�r�U�Y�C��*�R� 墤d;9������Jt�d�e������W�Cbl~��F��ed�R~�w<�s7���IZ�%�.��i���!���Vz������"=�A��ҵ��Ls�s�7�|�T;���bQ����x�쿡���3B���K�%�u+Zq	��Q=X�D���fD��]�� ���̮~�	 f��M�k\5�9wBM0u����O�c�b��QI���RJ+�,��$N�|pxEX�{�:�1�]�}�ϔRܸ�)_�h"9��wՐZ���@\��WF�:�i�|
8@RG	�������H����3���n{�j2�I���kZ��0P$�]��݈y����>��B/2z��h�|���kmǒօs�M�(�O���~���~�ęD?�~����HP�w{W�*�-�I�����D-�G5���i��]�{�/��r�HSW��r�踵��u��P�.�B�n6i+&m�a[�#0ZsZh�Q�Tr��s��Dɛ}`��ꄃ�����FB��&j�bg�1�����SE�þs�~)����%�=x�^	��������;K��`D�p�a:P�xJ�T
MC����5��%���/�qp�T�5�n�o}z���hmU�@�~3��u�������xg���\j(Y�����fYv�+�t�[�Z5к�\g���r���|�A�&�����R�^�?6���)"վʓ���,���|3�h��S/�p�Չ����s=��G���6 ���QG�dO��$�� ��;Gv#�苭c�}�q�pYI};�$�vY�Vo�V;�}ZV.	 ut����	������Ʒ�x�X��I@����>Dc�R���/xG�y�Q�f��ܦ�2g> ^]:�e�P|�; a0q���GD��ޚ�ZN�N���}��, �WZb�%^C�\�޶���2��1���ߡ��nq��Jyx��Mc�_�a�<��I<�lh�:���qȽ॓�,�{�٩��k�� ����|��Ψ�W��ُ�k�"�i>%tw!j�b�#/����50T�x3[�����yn����� ����~�W�5�&�L�ӗJ�3���D9d�Ȉ�����S�"p�4|�j���{�<���Y=�h5���
1(�rE����-¤]�� /�ZM4z����鞈�T��ޖ�����N���ҙ~T�#T6�E�/�'o��hܗ87T�š���n:�z=�yi�+Ӛ/��$�U�	��K#���Ko1��P~���'�	�#�/^���|&�|���P���:�h���ŭn�Y�S3rhu��J�y��]��k�թA�u.��n���T����q���G	�}�'��RЕĲ��&ԑDWvT�F�Er�b#�&^:�� �D`ۜ`;ۅ{ſ�n3]�7�X�X�{�{P�D�}M�a6��F���/�G�~��Y�BK�}�Q ɨi-_*H{�v�o��0J�.��y��ap�c�	&�oh��Ĝ�C�{�Ρe�[r�Y���Fԍ㟁��s�cd����.�T/w�J��j�9��AE|��V+�LJ��ܔ��-�$̶��d��矄 2^�Ջi? gx�{5��|n���4�=X�`[L�o�ŝ���Pp⧦�W<�ӎ��Ό��\'�q�;O���9q_Q3Z
�;� ���(������&~j�����}��6յ(L�m��k�=�A����6�n��1E����"���K�(�ܸ#K��T�ȗ�*���b��?�_�7����B���f����#R��Q�2^Q� �n*�P�,���i��'���2�,*c�c��Ō�.�6�r�I�kU#JA�R��n>�n1LA��-s�<���d�3m�u�t6 -�.Ԩ��ത��*/�9��$�$����f����L�x���;n�����rQ��2���5���*�7(!8�]W��柣C�[�ֳ��nyN;.h�	�,�W�gųF���b���!�?�.r��q��3q$l�h�-��s�@���>�r��I	"��l����Ǽ`��w��t��q,����o?H� �5��FjOn��0�)c��;�#r7?"Y＇
�G���p2���I-�P�=�Յ���楃�㻴�O�Z5�p�� ��A���Աw;��^��VT���lc��C<7m�/o�m���}�7�$��DKZS�o�N�@*4�@���W	s��U$��Wa;�=�2�Rcuӵ�����H-�l�Ȯ���v	{���`��m��N�Lb��K��Q������w;Q#3s�E�vzehm��s�ѥ����S,�Y��D����`В���͠��)�o;jS2��UgC�E	���y}b�z��a!/�(�4M���I�BV��٭�f\���^C��l^���n������P,�|'l��D�>tIe�_���_�-��K���G�źځ��<��k��hyZ��[U#�<�-B�/_�0 �KbV�5k��]B�"XV�g%�I�X�*�RJ]����Ӗ�� �r�+�����jO&OK	||��d���bLpFg��xa���0%u����=���s���u߰Qi௜�"+vV�)Lۢ$��p��À��)e��[��@%���	�eL-��*���������͟�;(Y��J�����Oz�ew�o��>�fj��ɋG�� ��9�Hĥ��t������bx"��7}�0kh"˄��/}��Z�0��"��������yU���:��̶$�y�2��9���N��˖l��Xߦ�C��2��S�(C3eܙP�8b���ح��j��chr 6�0@��E E+Ci�%:Aۗ�v�$� `/�㱂���ŋ#���Lb����@�8O��Ա]�1�I���ߴB��*��&����b4M:��w��q�8l* m����N���ҔTuA6 &�zw(��nV�,�`�}� /�Y^�pV����v�U1�q�|p.䝋��4��X+ZDE_m��F�`��w8��<�b���n'�O4KcZ��޺�S�8lA��O����r������
ݛ�,�n���+E,�0b`9"�� �KYT��%>��5�cژ���'J��X����E N�{K@a�jL���О�s�lE�̮	9���i+F�L:D[pH��SU��*M��uv��O�G	�}��x�OCE��.��#�+�Ԭ(e�@7R�\4��E��%�S����.֜P@*��7'ۢA|+W�w������H�;^���
촥i�َ��v0��֌��)w�ݯ$>v͓�/6Ru�3m]��A �:鐔?��b'�h�p��I�ԑ̫��u�� `�ka� Ÿ<��v�%?��	����N��X��n_��x��H Q�i\��R�(.�S��ڿ��[��/�Y�l�*�w0��
�[|�=���JB��?�t�� +A�_�M�\I�]�*;�Ѻ	 FCo�=�W�)��l�ْ֮���@�%w�n+:���;GR���(^��9�\���4)�F|{�ϫ�.�(��,'�z��!�
`P�T8�F�<̃(L�!\L稇ci�1������oH���20j�W�:�$C����4�V����"�%d�	���A�}��*%��m��g����m	����ݫx35���4\����%[(,7���fh)n?u!�8rQb6�SU�Ԥ�l�E?a������~��[g�!�Z�������ǒo��'�b�����L��g�-?)=�kK"s�g���,�1u� �h��wv+�W��)Q_�^��Q�����^��~�� ����	�1.����c�H2���Pf�[��C-�󋥣�,����C^���d��YH�<S��R�۝����[�_��_1(P@	t��:��)�Ȼ$�ۥElݵ5�������T���CtMu���6�G� �L9���N
���dG�<��Z�'	�ѭ���y��gh�^�,���T�H!2\H]����]o���rr��1J���s�ǀ#��X¶�������O�|�v&�Mtvw�tA��V�32-�2��6]�b���9ZMy�M�ϸ�;��S�~��N�Ź0w�'Ñ�6?�|�W��K�#�[�y2
��h�09V38�K��