XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���<'aw/�v����m�2�
�ȗ�,�H�}H76� ��e�fF��~GqJ���qԡX
����M`CY�Ͳ< `��'�qـ�F'��s�x?�:�γ��\���������2�.�f<|����u�?O��/ȉ�l�KV�L�UhU�w�k~��M]I�$�Y�ּԧ:yF�'�m�\~�{�:ړ����3YP��GK�����ּR��pz�i�1b�����7���\&+?S�3�1��1�Wte� �����"8���KI�u ��T���-�8�6� [��z	Ak2ZX)P��g��ۥ��+0�m�k<W���.�
mx�O�Ƕ���͘�
�^��Cd��B�o�N�mT�����EskʏȞ������^n��]nu[����׀�S�5'�+���|�����Yc�����^/<�E��S���S�o¢Uw�5־lwx f-(C��)�C�e���O�	�Ӝg��}��V �L��z��!��[�F6ղ�%���1�!���҂;�|'�=�Q�U���"�ꬻ��a�:t 2�����(�Cz�ac�o�˯�)�ޕ61�L�p?�ԝd�	�au�>�kE��a1;��cf�ɂ;5j�K$y�t��kp$O�T�s��HU�&����(�)*0����
:��m-6�"[������@�n�:���7�^w�f�9�� Kӄ�z���}c�]�6�&���֭�͠�`tn.�A����1�軎��wmx�1���BXlxVHYEB    8388    1740^�st�_;@�Ű���ҳC�z؇�T�'��[����{$���P
�+5~R�?�}�4�	����L�����*�sIz�dZo�"�:���<MM�=8�q�.R�շ��[��q�Z4��+�� ��[�>��'�g
kO#��x�ҷ��uҺf��R�Ҩ0V�߫~A��?�jM�5�E�C�nT
9��{ӷ�?U)�{Li�7��BV�P� ]6��4�7���a .��dE�G%͐L�2`��&�E�	���x|�6E1;JD#:�ؾvA�9w�M� ,�O�4����=�u� *��Ͳ��33 p4�Gi�C�|Q���޴TD��	��:�2���8v6F��$w�w lc�X�Ge�ܣ�L�-	�ԢDCn3'#�db��Q�z&��Q<�ܒQЃ����V�Ď ��?�-��ңc�KG���T���u��p�l�/'rw�La�-3�����-*�C�*25_�5+� u$����$恠Hj����UR��I�2�7��,r��5f�2�ɜ�I|C����~,m�a�JX�6kً��>fU��l�*��삐��(-�_#ʂVw&E��P�F[�N�l�91ೢO'�C��T����Ad(v���f�
��3:�	P��1��wRts�.����X�*U��=�[��a
���)����z�x�=��N|u�[������NK>���� ��5y�]�J�O�c��;I��ä�{���d�6|6]��Xn'�_E��Gw���55|�����j�0��u� �nA����c�(%�K~܌���Eo���S ���N֫����=��|&��#g_���rS���u��v�1��O��3��O��w�Y;/+�C�I
����w���z��ħ����0>}�{2a_�: Q�݂�5�Aoi���>�83�`[*�N��� �������ؽO�X��m빢
|�#�C����7��J��Ix�`�lP��UW�0{�{�1ɣ��M�%�b�>(qk+����h��&�-�.��N#��)3�զa�7�T��U�l����&������r�����B����<*"5���.�ku��S��|B5�!�Vs���m�n�n�w��}�豾�5od��=��a���]>+�Z2wVgcj(�3.�Ag���	��P,͎��?i�;�ޯ�y�[�`�Iz1>;k�8�;��i��?���Qx��j�c«�b#�]13됑�	�^H�(^�jB��꾼'�E���W�t�g1������r:��D��H�ɗ�eC�l�,ߕ#�#n�ʹ ��]�g��N�)�C�;��'s<�G�5{$B[��ה���M�d��Ջ?�����D���mlu#�K�hGD(
b��7@���Q��o�g;6��n3�On��KO�wJʹ�=��(�����%x��	
Ձ�h��/[e���E���f%�X�f�~�Fy���Nv�]Ў��d'q
PK^�z�X�4m�zb������s+�ĝDfHHB�R��ժ��m�ry��[;~����+�L9}ZJ2N�s�$��EQ�%��nX���Bj]H�Cn�^M������l�=�`�Q�	�o�������5���}�0�x�Dg�G��4��S���ߛ�Gxƅ`C���m	�k��L�1����� k�s���խo��Ͷo8�6��z��Uo $�Y[�@Q�)�>;OŐw`�`KI��Rw��9`��1�l��>�U��=���_N!��bh���;��>ӟA�Jb�To}C��S�^*R��G �?@j��3,��3�b�NPEƻ�%4����0_7W' �����Rtoc�~��j̍��61�54/�}�]� ��v<�>�/n�at����q-�� �t���ˉ�#���u�c�L�obȍ�６ i�x+���vpب�UDև�o�?ZB�y���T.�1|�utj���Kث󦻤�9g�Uin�b-����F��Q9�ȩZ�2M0�����l��l��=cK���b���OM��@�!m�*ik��:�����9��4*�]|�u2/B���"+Cq?U
%���R�z�!��WOiF�YV���@C��E�oef�6��b�%�|��3v'����st<�"-�h<�I��̓�
M��ѩ4��J`��m
�����������6z����3�{TJV��R��1�r���������T)v9Y�����I���q�0��ۯ�&s�|��<gv�~�����I�1�Ӝ�	X�ؤT"BLs��|���z8̭�5A��狃�o���o[j�j�$�)!}�q�-���KN=�۲�>Aߧ����Z77���^�{"�PY2-S2h��i�S���߀�����<@m��M�<"���c���vZğȜ�<Y�T��5K/�s ���q�
��4�_�b��BW{/�����S߁wT����ϐ{����ȳ�X�5��M�}+�--H_�W�T¼,u#)�o7N��ak`���I�P��/��u���fR��y���V����f���gDn� 	90�+442b[�*_�T�rCl����=s7���M�Haֹ=	��+�� ��-b��� �:eW��� c�����4��Ը��O:E��G"��g��I�O�nV͟�uh�T]�0��3w���$+�-��BQ�nK�N����^T�Ct!fc*"���x�ɷV4��-�˯���jӆ^&OX<S�kݵ��r�G�3�>m���&�ɩJ)eXc�­��V'Ф${�����:�En��9=�T�[�tT����P8�ͻ�.ɬ�gs�G�#�A/�&�זH�~�*�5���9i	���e0NgF�X�l\"�Ag��<�#A�G���N�*O����B�!t[��Y��H<��_��`�o��*�%#��F��b�����M���x�A�ҹU}[n��-�w�KZ��!;"ӎ��u��<�U��y��xQ����5��8�o�`�a��Pq?���H�hZn_��>Fc=}ثA&=T_3�?�<�Z�ԭ��K,��Qα���ȫ/�ۭ�p�ˡG!��0O�mɩ|(=��	�ǩ��6=��ȧ��$#�肴�Ml*5i��V�σFߴ���HW>��3^��3�&�۸� ;q)C4�hB�/���^��6vd���P1x�8�$�y&�kN<D�L��c���{�̠>�	�P�Ch��i�`d�6�li�qfq��E��AV螦��� Mo�z!Y?�W�:N�D\B���һ���/��;e�B����E������@:���w��E�	T\Y*�8G��I��@�#�K����r#&X&�ܔ�����yŮ�����؞7b��=�R�`�Y���"��M���:h�2�V5I�	��H����PRycy�G%�o��,_D&|&�>-�0�>��)�^����t�N�uh��T)PL�9CT���.��Wɹ�����t_/(w06z���@LM���wbI�F1�dV��}��e��M����s�dt�Ͳ3��������π7u�u
��^�~��n�?��Ho�<�
h��h���*/g�5����sۄ�=!/��P��֒�x��r1��@���Q?(���ȸ9���{�����P.��* O�V��?�0�3�n�rh�[M	DaW�' �3�}HP��\C�[Aq迾6bǤ�(�"t~�ZfD����,�r��q�����V:��t&����u:d#=�i��R)�����B��Ḭ����
#t�lp1�!E�K�'���ӡ�����g&sU��gs2��|O�9�S/C�3�(�x�Y��@�>0���T�#��5)
��6��	ڿ����@?G#gK��'��!gͨǐ�F39��������ԇ٥s��U�����<�\yL|6��츯ꨱ�k�;/_jE:y��R��۹Z������L`�gtT%�����ɀ4�"��p��N�C�j �B`�>"�J^=߸�1��Q��V������zK�X�2�x��&8�Bm��tu8�E��Ɩm?�)�r�gv�o|އ����e�W/�ҲH�������S5*!S�"��[�_��i�SB�/�]��m$�*l��59��rfØ�ž<�W�s)����"_�DCਟ!b�l!�
�B84I�<.�I��K֔�34��T:�-\��B`����p��K��3�C5~�'z��uMo�����(0j~��+RI8b����B�"��v����6��ރ�J�ʡ���A��|j����G�
���1{ƾ�(������g�
\�9��Uwt� !��x���6SӍRǸ:�l҃D��SR�0=���x:$��7�D���[���X�@4�~~.X�y�������&�ߦ��.M�R��۽7y����T6������:�W9�"������԰P�����T��|�S�I�U�bp�D����F��Z|;Y�0?�ʐM��6��7rc�"�u\��nQz�[(?@�n��5nOHp�U!Q���v�:�����2�e�.�	C�8�+T�F2F�a�O��c��$�1��9�
�}��q.��ER{$DF�@�'��<H��g��.�;�����t-��;�q&��eT���Ko��R�bT<!��κ��c;�!����-�eo��n)�n���F@ƒQF�'�֯���`����mY��l�C��ik�PZ|���
��b}~W@$�k�}ϛg6�|G�8e�Lh&B�x�d�([\�薎h�l��µl��TE��/^9(2]�2�7��$S\q  �~R-�����+�ī��@�X���]Q0���,�f׭����4��M/L�Bp���1�+g��4֡P��j���bE��\�@ѠQ�1~�ܫ���=������ӊ���6^�z��.@��ԥǠ7��Q�,B�.����]���8%ؕ3+�і�<����"����#��3���`9?��z�G��+^$S�ip�D��=�Jr,ԁ�QYcJe tB����g,�q��,�RdV�6t�R�2�t7S�5(�n}��M���p�$���#$��$�i�nX/�L��B�e�מ�ynO+Ծ��*�� ��o�ȕ�)��x8����۲����1F���C �]�?��'9�*=P��sd+���*�� �2~��m��>��lN ��x$֧)GЍ ;0��āA�
��4/��-����
�L��j��CK�^ɹ�� }R��|�bN��͟��ߋ]����zmn	�����ׂ	�Y	���������X�1�-r��H����Tm��\�!��#%�8U���H`�q0y�۽�I�h�P�(�4*��S<>��]��p��ב.z鯯����_�8���q"9�x�8���脴@U�ðDPh���N 2c�
�,����p�n��j��[!c�Oe@�K FKc��-^�F��H	����0�l�J�]�����*V�:�B��<=�x
�1h)��E��@���e�Q1��d����.�;:Xm�r�,2��33a�����c}
�D�"��Ѩ�l�cQe�u`ˤ��"�K\�P���yH!}�x��/��j`�R��-+��$�*dV��S,�a��Z��urY��,��Ѩ�wT�s�X[��;�K؇�X�Ncy9��J~Z��I ��4/ʶq��x����d�#Y�X���_�����(��E|��ӯr�]!�}���`����u`�(*՞6G�D���B;I{��_K���D��@����-*�\����&��/������V,�cO.%_7�?�f��V�G�=L3�ײ/�\1#��?�:Ė��R��N�c�c/{�mn��.���B�N4S�D�.u�w�w%i$^��=0��֡����