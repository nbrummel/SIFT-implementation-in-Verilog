XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V�����n8�0����rL�َ��F��țZ>4؛ίǣ��/r�z�bzZ�K��h��&ªc.>fl����	�B>���Fͮ3�H�)��bκzU�ef<�t$�C�zC�7a�`���{b�,C����8��p�,����^�\�"͒ �Ҙ�G�����x���ҡ{z��F j��T�dʥ��8�@'���6?�07!*$Ά��9::N�~ 7$I=���8@�鵄G�X�ܨ���X��@��O��`�+���D�PP�Ϩ�=X�w���|8>a�pX��'�j���}�4��-p�B��q��g����X��6��m`�}X!-�u�WYZ��-Q,b�@݊P����ցgFGg!�-=d,;t��˩QԢ�Ou��,H�%ko^^�}8Tz��S��M���Q��J��'��g��mN�r��k��IQ�I>OQW�Ǘ���j�1Ʉ��O�kH;�kICKOc@3����+��������vz�j�ga`Q��\>z�`��G8�,Y�e��Z���Wm'b鶇D���5"�'e*��aw�)��xb� I���w��=��K;$���E=���d_5ؖ	@r��֖�ktƸG�	��؅��mU*LV���|�3%r�A�gn����� F�Oy֖�Is|�`��FQ'Y��j�xF�W���ߝ��'�b�w�zj�e�`�MnS�f�n�A���R�W�"�_�	�y��Z門EC��g���>PV��r��T�-L?�T���d������q�i�:�$q�XlxVHYEB    c3e8    1d20�����n�_��-���'�`jޑ���������!>�ΑB�G����w�SZx�ԇ$�)v�L�<>����i�����v��]|3����t*e��՝]/E�,iX�B��C@�9U�v���8������i]g6|?��l�"u�
ҟr�ݲ�bn��WH�j��;# ��<���	��/߄.������ �A�n|��	���B�3�'vX�����2X)5Wkn��滥r�Tw�g�s����V�'$}S��s���a��C�d�@���}*]zwj̉f��?��b1�g����>�� r�w�7E�.�G�[ʿiP(���Q��>x��`A��ub�?�������3㒳?ff��Z�	a�;b���n@]�Ca/g�^���-�T��IwPF��Ci̤���N�͗8�U�V?<�ij}��Y����������(O��y�o��z��gzhm4����E��2U-2�����$�FϿ����G��Q��f�A\��9����mr�?Ny��@W���R]�l\2v�F�6X�����؊���+�^9A�
>s���M��;e�h#�.�l-{���qu�nlJ��n�ݼ�o��`�e�ii��U��<R��F��(�͎Z�BЏ;���Ό�q�����N�v����28Dh�0qQ��+�pZ��P���.O�������_�w�Z���GX����%#�=WZ���<a�8C幙���������l~���Q�,5Ar1�Ц~��)B��Tm1d�z/�����uO#�vX���f!6����ǀ�����45���:� ��^3ͺfQ��M0K"]�~й�����#��O�O������E��)p�\��R�!k��w�s����ŋ?�$�o��p'�lv���F���nh"b+��,���2h8��^�+�C��t0�P�ĖбL�];��ů�˃D��<=�-�������%�TUet"8���o{ ,��LEV|���~M�id@0�ORم�k������q���)j�Nӹ�6P�џ��(4�9���$���s�"��9������񅋵dlҩ��w�%[�?���.-��ϳ�����Ww�e,������2`��Z[h�*.��>L$�?G4k�m����F�ߎ8]�b�e�0��Pm��V�ύpcf}��j�	�Շ8�rn�D�����ީ�|O>�S�;]�4�)z[��x^���U�lmfX�o�uSdh��[\N�q���ؕFZ�w���<��SyQB�.>Q��@X¿ĕj �֋�t�� 	��>��-�R��{q���CҊ<ݏ��YSK��>Jпﵚl�Z����\��rd*���f��cow�)��&��k� �c�E����^vVF�y�m-f�(����hѴ�*�Όl7�Y���K�1_��YM�

|��pFV#�s�vD&4]��P�_r�cD���<�?�i1'�w*>.���7�AEq!�O5�-M;K�%�����g�oZ��7��;�"�(�m�� 0Ϙ������D3��Y֧\b ���fb��IZ_���ӻ���J�?,�KV>���L��8o��7�����X܌pMn�7���w�p;u$�W_�wJ�����t4�vm�`�W�F���Ո�v�dK/��|�m���$/�6�H�g��w�.�E${x�3䝕D�g=��پA�aA�Rȉ[M�p%�V���_~ܼ�ں��^.��_��9���(�$l�2���2��������9������D���YPa|a�`Q�#���V��v����>1���e��E��gӍ�U��n%v�E�7֔+�e6�c���.����9sE�{��3b�<8UmJ�gA��ߺ;`�;�M�Lrj+c��^y����|K���:�	?雔@p��ͧ��i��˩�3{�GWr>V��ok�Qm��%u�ŀq�jj�
��l�`=����8�X�C�B]�
������=8��fi�n�	H��=�I�B*I�����ط�̈́A�R@��|ge�AM��n��e)�(���sM��@D�3�j���?�m�I�Fv@�]��L���q�O�ڐ'?a�9�i
� �T�9Ey7a3%9ɮ���]n'�w�bȢ��ɓ�&��Y�� Xm)=J� �q$�޲�<5�:�[ �t,�J���/�` A=���5'���O{�\V�x-��O�𡀓�� �D�1<�fX�j�L�z��曂/l'5�KXt��2Yn9z�5���g��*Y��@v?b���ԝل��3�wx��>i�����ݱ�.�"F=OQ�+��y�������-nDg�<ģ�x���,�p�5�ipu���H,F2g`U��;<8������e����h�ui�����E��/�a�ľ�{H.|� �]h�	,�"ل����i��>�3��K!��d;����ɑ�
E��+&�i���C�x��@��\���<1�f��u"�'���W/H§��-���EL6�l@�Y��H~X�r�4�%+݋�1�[g��J����G�xt�� ���S2=��WY�'9˲~����*��3�CT�ǆ�1D?\ʖw�q�9j\B��e��G�愝�.낝eԭ�-����{��2]p�=�)x4>I��>��y`T���wQ�z�U��	��u~�Gp���z��	i�ۊ.٣J���(�j�&�$��TU�	��:Q�ţI��Ǥ�&�ǀ�B��t�a�b�c���XPn��_�~m�D��KN��R��x @H��E.���@�{�Ï��']w�{��J��:�E�%�%��+�0	R�A�Z�����u���^v����2-���rh%;��ǟ�1���Vк��a,���VX�ۜu�Wʯ���� g�9�Ї ׿-50��ِ��rG�|���y���$��{P�r��)�91�����O��O��j�'`�x��7���zO>4 �-�����Ji���t�Xg�����k=���R����=u�g�}�݆���q�h��D��$6Vr"�{�,!;��3	�a��y -��%z]� �}���2�A����pSh`��|�}�㑈�"e�=��o���#~5{��c�c��SY�/I���dM���cU��щ)�s��d��f�����?��hIX�2	Al��怞�[�
9[^9��4)z���<��Ȼ�j�l!�=�T�:�a���t���&a��?�O�C��X-�B>'�9|6Y��]_��RK�p;�꾗L�`�� s]�N��}ZO�������	O�~��5fG>�ɢO^]�~L��v��݉�8D$Ǜ�)���� 3ˍ�(�jnq�S�ƽ�vZyg����p��5���NM��맜��U��L����b�U���޼�me�H9غ��3W'������#'��ȱ�#�W/���j�;,�i���p~� �j9���t�`�8��*]%ɹFP3�����N��rOg,�
�8��P��ӕMxӇnb6�ޠ�è�m������ؘu��Ѭ����"�f��K� `F�|)�cή�e��-��D���yg�/jHKeHr�j��p��tR��������o��wHD��bɽ��9�3 >B�A�녽�����y�(A����\܉
Ԣ{�Gˁ�w��o'�W��.�Spc0�|*��l�ǔ�$�M�i�i�Co�� �8���ԚCU��w
K�+��ŕ\��]�Ȋ:5��Bhv~|5��":L�Ј))�Ҧ��8�ԎA��8���}���(pkf�(�o����>9>>�qw,�0�2 ��4;�;}�g�NP��-����mBaDDDf�N��;>X�8Mr ;ox�M'Z�w�^w�s�LRG`B����@=ާX�|�u��H��<S�t�HI�r�𰮔�S#��vD�p��9�I��e&���\�r�}���_���O�\��F]�!����,!�q!yV�<	�j�bZ��@"��˹���9Z�J��'�As��x��� �h�n��73���3S��=^:F#M�Y%{�ji�.�P��'�	����q�[*B&�&�
�\x�\I�{!haf�?��K��H�蝴���ܦA9��ۊ9��:��Za���ރBł�NT�<�Ύr
�mO��,����9*h��;�����d��\+��ȎV)�/5������@���\�ߔ�"�|P������:�Ea�Q�.M�IU���{��&��!����۝�[��У[t2p
�lG�'1���S��_���m7�@�%laRƛ��+��#k�7���Gr&_1�%N�Y���9Dr4}$���i)Y��/����m�tp �݋�	�T9����"�o���I���z��
�����rp�
;
:��x��	��_b�]6>�  ��',FF�T���| A� ��J�IF��2���"�̳f�T��_�<fK.�R��#���PGLBӡr�_����H�o�U��\��-GH�R9We���: '�N$��+�Ҁ|�0��R���	�u���2&Z3�u]��;[yf�1hVnȅbn<��iأ]*�lؖޔ�8�B��8�@?�������>��dǉo9�(��f�J�bw1���u@:G��H��'�7�FPf����}"I��&z��5,ey7��SJo?�
����>��l���g8�<�H�ޢKZv[��0�&��`ˤc=w�T��T(|�}���/!�.�Ä�W�:+��~5�� �m�"I��ڃ���ّ}���g�H?�xq���EEU'��0\lrJ74����P���>F!k��;��L��P�v��j�c��C4sy�u?_��o%[��e��L�Y��I�����l���G<۪z\.�YGƫȡxl~V[�j��dG��ռ~#i^��~%�቗ze*��4{d��!�6C۔b���=�ُ�� ǙT����;�̿��{/�MG���]�K w������"䦯Z�!G��� �SZN���-��`*yZ5e�6�W��.�㮌��������v���{�����i�m�CԙL@�V�O�;�w�G?�p�W�V�Mĕ�sѶ�[Z���6-�&2���'�� x.��z��,%�t?�����b/��m�-��$�ެ�):L�����:�o5ו1�t]� ]�#�s�=:��.78���W��~��ۛ;]>�~RT��f�#Ӳ4)�9�*=W��J�s�ȫ懷�>��B�ari)�R���U�4P Ѐ�6f��+� ��]#g���/}�	3{C���[����cw)�Z�(��f����v�3�|�"�O�Oy�&���Dm��𢏲��l��$B;��9�΢,/d	�ko��Q�)p��m��:TYC^��.�]V�r���+yl����|% ��j�����Us����%e����
ot�#�XÂ�����(O�����0�gw�?d�HVy�z�Vd��F�|)U���J�R�f�6��5����Gy���׉	!�RZWy�l��[��؋J�)�f~/?��e?)QM��U�jjL�dbN��־�<&�K��|��=R�	��Zr�ݵ��*[d3m	Ƽ倪�vo��P���?�W̟����SrpN�L�������I�-'�j��3z�h~��������?���c��=�|�v�-s�v@>V����ڔգ���~��i��N�����3�3"�J5"IC��^��kS�y��bN�)�~����w�����.%����qʾU�SP���ΌU�	L��u�oμҪ�zCɲ���$ݘu�����4���]��D�3j�g�
֩G�@X�w��9)��i���)���~D�-�BH�s���-[n��|��2��G��'K�PHU�I���`b�s�����#p�i�X���2�E��+�]�R �E��* ��;�W����i�R��T�.px1ߚ�QN]^��i��(��yD�a��K���(B�]��Pa��J"��~�v�/L���k������*�@9@��0�z��8��@��9�
�舴�@���+(���Dfϼ��	tX�8�vG�'���A�n1�AubT,�J��I����U��C;D�I���֦H:}�j�` v�EH]1(!vl�ʉf�d.��*۲���#���e8m���c�u�ޥ�J���l"0ۨ��Q{?��&(�Q��J�giT�T�&T`��0�ۅڞ�T��n#)�|��m�Y�.`��nM7"���s�@^�
o����!J�F)$4pU�����^�1���Ęp����SS�׬J��1�)x���g��C��-�b��B�k}���s/��S���񭮂���S��\�_��֟�바gR=��IZj��
��	�h`��j�B�Z�K�8�@�����^���9�j2�|���������c]�.�Ǿ��?�K}�sm�'G���ՂPF���R]b]��=� ����L{�DԾ��ive1I,u��3x��X�f�FWI$j�y�'3�d{���	�;�$(Ԭ�@~kP�.���,�*)�^��vt��ޕ�-��1�=�jS���@��1}��㴭Y�qB�z�J0�,���j�ޙg�
�q�ƪ�^_�Ί(֛�Zެ�ȅ�O�ޅ���f|Q�_<��a�B3����(fP����a�2h���F5�<�h���0���pt|-��N�z�G���$4�_NK�h�PKS`_9���~�HEb:���b,K��+������I�kJH4�I�ԫ��;�(Yv��Ô��Ԛ�G�59B1�Ɂ�^����?�YO������������ڣ��S^-) �)7��ٕ�G��C�uc
�����s�����}* {^卮Um��6Z��-!�4 �~WG;��K�<�ݓ��Y�������`��NȐj0��+��:O3�J��]�s�]���'��(�&�o����X�,[ ����vH����]�?t�M�u �UUr�.6�����w
%�X7����Kxv��/���wqd�_Ǝ�)�2�5QƄ���Ԃ���8�;��W1���#��A.�p��D�\��Ljjg����@���O�d:����A_o4�X�{��p�aHD5DHS@���B�j�˺�2{k���o����/����Ul�:��)��a�XV�1$:�W�|�:A"(a_{[g�S���&ޣQoY\�'�g�b봅wf�:nn8�3�B�G��O4��X���Rq���U�آװ�����y_������b ��7�x�����sA�E�a�8L�*�sɖ>ċ��0��8(RS��R����k�;����8F3����j�ﲚ�S2�ԡб^C5����Msc����Q��