XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/��怡6�/����G��F�g��I�>k�^|��Z�3������e�~�G'~�< i��7�o�+3���[�2�ym��>��d;0;e�V;Zd��c�-��������7b!F��r�������u����ҫ�n��C�_w�p������6��J�7:�N�/�7�g������D��
�&������g+�.�B;ٞ�.*��t�],�yי|)�F�q��~L�M�톔�'̺�Z(Z���b�-��e�0�j�/��H�/UɾH����c����~n�|ZZBG�0��$�����_�����Ѩ�O�)g�4>S�9�o%��y�����m����4�܂��m�Z�$�Id�p8?�Ont\�t^��I��"Z��b��� рK�;�`�m5B�ޱ��:2TA�"��E8�fxs����>Ut$�b�1y?��UY4���2�W<#�������Y�iB҂_����7Fc9-�+XW�ㄞ�q,�ri��%l��?�ea%�[p)�sR7$��0���W֋vϻ�a�~�"�x��N9#	���o��q�U��%����Eg�8��*`�ԣ|�	�b��8ORt��mf��e2��j~�!�O1�Ċ�<j�l/��Qo@�^���W�U;I�I/<�`δ]��g�s�q��{��ת�7��2]����
gQ1��/_�ӧ��)]K	M�ͼj|����+�
�*���~���b8�Ux�V߬�,��|�_KOn�ExD�]�� �1A����f�蠂Z�D�kXlxVHYEB    1e9e     910�~��oJ슰�Ϯ�v�?��΍9�z#��B�0��6�.��Ya���eJ@>PK�t!�j�`������)ҏxu�ۻ�z�u �_c*�Z�?��,��q��J�����E��!>�e|dѿj�tuSl78]��[�D�E�� ���!�����F�%n[����������Qz|����;�xJ��Ed�DQN�[��ݡM��MuE�Użr|�� s�!y7�W��&D�Bo!�41�Wv3O��d*n�r�����G'��gV�x�b_�5�'�"@�c��Ͼ,�Q$W�N���3Q���&?e��D�a�b�$�ihZ��������[1(�P��Vا9̒���o�K�G��.�j���Y�}m
W��n��n���@�F�6w>`�?n�yL�����YX� ���|� Y��>�0*�q��q�K�@r�~��1_%L�E�Y	<לm�&Ĝ���2����ō^�Ө9oN�����I�
k��o� �Z�Q���}�٦�R�=�<� ,H�@{O]�*ĎX����Yyƚ�jSH�jyI����l^���&M%�y���@#�����-����dd�xP�C^��ҷ�4��.�;����/�����6�C���C��塣`��_
Uծ�sр4��b�O�]��@9�i�G�mw1�Ÿ��k1 �0\˺�&Y��,θf�1ʨ�u~!n��\M$&ͪ��ZP��M�.���1Ho�t��p36�7��@�>��X��&�Y/5�H����_�E��r�Z��Kh���ǧ������$c����Z��#��C^�w=p8�|r�5io��}Aޮ��F�����X�<���Y�YK��1�e)�0����@8����6����� �$���q
;�Jr_�%�1\e�|�xa%���LZT�,ne��2�?T(�p�D@��O	�3n��Smb䲥���Nd�����"8�*�3Bӑa�sV�[X���_w�"�&r�b��ms ��~ �_��]j��=�I
[��gY���ʙ5`t���n��g�֤�'t�Q$G�]�%�3��f�m� �� ����ہ%M?�:�c�|�&�k�!�?�.Ig;�T[c������AS759�H7?�JA%�H�T�]�)a}��S5v�]�_�6�����\�s�?ÃS��/��v�/��2��M��̈J[7v����f�v-�@�v��F�WS�͠c�a
�%�F��^�6[��S�b�9��}��T'.Kv����o!�'����)�����jCTM�ܼ���wK؈e��=w��WVq�4Nz�e4�- �*p#=t�_PhAc����֎�}{n!���+�	�d��\�������
�E-/B�Z��#�{]5�wV�'�(.�m�Z=�`~�-�|��B�.`���!b���U~P��*�k��!_��9f�=�\�C	�"�:�x
������;�N/���ozb~/��Pz��0�л�ʛ;�mA+�>F	��5^� ̤+"�i�-�s_��D�|l�ʝ�+Aj�	,�i�2��`�X��&�]��=gD���xV�%t�P�CwݼKCF3n�{�͓�:��S�/l�"�,�ֵ�b�U����RcC�>8/�!�z��(�|���,4�M Z
��)�YJf$|`*K"ݙ�,}RwY�b�W`�Ҁ:�^�2��|	~B(E����0�Aˀ�[w.���a�����M�J��� �S��OsuT����Y j|+B�-o��ڿq���_��.�.,~~��g����d����7�8�?$d���B��	�$��=Q��:���uq���s͋� &�S��sݖ��渧#���0�yh�� ��몸d�6H���XZ�']d|(�B2u�;t��׋#����N�sY�����0Ć�oSͧT��|����%�m�!MH,i��H�Ѓ1�^���t�ڀpPQS%��y�fy�18��΂����ӕz[�v���G�����%z����~G�Ԅ���p+����`�����6�]��_3��_}/�_�G����^2���V��L�$��*5$7�ȧ�
��*�#�!*��C��n�X_���x��]�X��"xl�~�e�A�0�0>c7�D%�b�o=�t>id=qהNa��ߊ����#�+?� �ؖj�$�;�����<�y����OzY�\tB!�5v�����n�� QNGǽ�j��kkb�����WsO|��J�H�7E����놻��b�5���T�ޢ�hw�����w��#�l�ӹ�/��:Z��