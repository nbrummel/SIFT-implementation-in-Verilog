XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Jw�����D(�a��v�T���G��$��#���ٓ�ʙ;�p����Iz���2�fa�"��TPW(��P�����s�����;}pG�E/���@�V ��t�����{���@�v��3Uh��4l��1��\
\f�)u�z����P�+��;w��x2��҄���ofB��#�+��Rw{ ��XY��ߜxb�^�|��ļ͎�/�<��h>|�v띓71�����C{�d6�Nb�ꤿD�G��*j[��
,�TF����?�5�~�;q�{ا�w��6�%sO�3J�D.�s�T���R����(ؓ]���*p�&��;���6maGיuz�Ŋ������M\N?�H�7F����Ξ:�@
v>�7��W��uݐ��n�� 3��{6�w�<��7�R^�w�D��:�E����=� ���B.C�1��(�Ը��:�1J���\%կN4f��K����W_����t>��z6�ٻ�G�:������t�Ɨ=tmT���d��L�,�ݝys����n�f�2��H\�`I!@a��o+�'�{�Ʌ��䥇(�0'��$���t�����f��^c��U�7����L���oԻ�]1l�p�:�(�h3���F��[\�"w"V=��6���{�@����(T:�{��?�^�����ނ�.�)K��]~}�R�i���gr�]zˋ+m�����p����߂�n�d���H�	6�Ҽ�Q/R��;��V�W���1�9��@�J���JC�3�OXlxVHYEB    1da6     940	��-ϗ~���=/�8�`@���<��a�Q���)���(d\lt��%�Y.���VY��8?�3�E#BK�
�K�Mŵn竐s�+r"+��>t]�(3Ow���k��Z�:��*\N�f���D�JFFS�_�z�{7�S�V2 u��Q�r���z=��V��j�W+����^���$D�A�2�eOl��>agb�D�����t �?���#�n�_�ugS\�~�QO^�r�ly�:}�l����^����Cy�H�S�����j�[�z[����ڐ�6ql:��*���i��0�L��ջ|�]
�u��H�rOEex���琙}D��#k�#ß��فҫ��j�(@��xI��b��s��=MFdZ�d��h��b�%,S���E�0#����>\5+��p:��6�#Ɨـ�!��������j�f�q嗷J��ܑs�6]ҭ�"��.Nz&�3�74�y�(җ�Pp�U����OdT� yTӭu?ʏ��T��.��W���p�S���,��~��?Ģ���^������Ηȗ-\<���*)yzƀL]PX�b4��Bė�kno�X?a��ٿ�^:��=�nʴ����|��s:���E E7���م�����<��q�=��\,��P���������R|��hw|���=��辕�����!�Kʚ��h�.��V�?b#[����?	���&��^�Qy��&B9Dy��b���cxZ�v�ꪛ���Gj��u�%����?"��߇`�:N��B�ı�xw��p�������=�.J}��E�;��8����s��zM�B�/:��JT\�����jAe�
�u�m�DG�$	E��TV%�_ �g��L���l,�)[կ�OR<f�>{�}֥\w�r�D��s;���h@��mlh������!��Mx���W	)���2�h��Ic�<$���=�{�}=*oW��]���b�~��mq��ߐ��Usc�i�KW�<h�o���LPt	��L��<J�q����1R��|R�c������=d���.�l����P��m��Уd�F8�_;�>َ�Yj<��QN?'�g:�*��h�,�W�"n���_�(�O��2h��BÅoA�QR�'���ѝ��pκe/�=sex��%Sp��X�}*�A��pHc�Ϲ�:@���)$�DМ�b(EѻS�m��'��~��i�h:�s
2S�$��Ճ@��_8�a2�	o�EZ��ȍUH�Ṫ�,��]�Fd�Xı:�_ã�0v�Qh[��%��s��؇m55�L
�2>~���zc�G����P�Δ=���F�J��w��+h�%�4BO�*M����th/j��������z�*~P�N�'�K|U	���V1Q�_�=��Һĵ�wX�DoA4��BS1�D�#x:g�J�/c��o�k�0�r��`C${P�R�2����/��Yqao��b����z<x�"�i�.��Ʀ��%��#��P"(�`'����3H�?��N�tٓ��{k,Lw.I�-pocV��0�`�����g����~G��A�!��wԌ�� �n�!�u+^F]��6E�7��уt�}ǎ�*�Nr�B�d� �k�˚���}����'SR��,G�5g{�7��q�4+��e����e5Ԃ�݈�꿥\^P"������8��'F��V�K'j�_Ļ;���c}W�Ck��q�j����I��y-� &+�u���1���p�"zr��Jfұ�m�g��$��=���Se���|~�������I��8/g/�澓�_�u��8�w�ݕ`�WQle���I<՘x�)�א_-�:Z��	����Ũje�=	�i��F"$w�
�b�5ʱ��T���t��#��?.��Q����,��/�g,A��rve�_��U�t�68�Dđ��!�z7�>l�i1ѵ�Jͺ�D�6�Y^���D[��t����ا��ɶ��.?Hd��ץV�06�7-XzcX�����C(
�;��B#�2��W�G,���D2�X��4�*�laO�t�扁����ƿ�H�<Z���4R��]���
e�y/�I����q��GȬ?	�h*̅�6t�1�k<�:u섾>�V� *��ĳ ]6N��>oT��.`nΡ8����d� �Bhk)P��+�r����d����"m�8��������	���VOn\�G��D�p��iw8_�u���4OZ����6�%V�Y��i54�%�F_�l�'�X���C�A����O%C)/B{�,F��s�4b���oP#eC	;���Mrb��@;��U����ڬ4��>��}�	��ԍ�