XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Z٩K�P�9���Bm2���mą=PL8C��X̅��ו�DTڽ/�z����XSd^=7���W��^��(����^�I�iK��:��'�ip���������3%q��A�trKf�<��^[֣��.iW����)Z�ȑ_z�΀��	5V�˲���Izx��*1�e�5�aߟ�d��l�7�����Pµ���'`]Wv��P>��5������J,��2��S�x��F����"���p��� R!E3
h�Z�7w�=��O,2��>�KW��d�$DO[g���됆��u���K��L��5bj����~cF��:�*B���s�L¿P̲�ۦnm~�I����ݼ(�L�"��$ʑ��U�����/CI���c�F+�j��:�lUx��<����9���h�`ha�ju�d�a�!�6�7�E��U��}�o$b-��
���!���B�1��8vղjD�4���_@ku��d�_�e:Ys�ݘL�e���?a�]��ޔ]�u+r�7bw��0�yA���FF�[R
�	�2<����i,������w�n߁w�>��s�Џ�~�a��Lx������/0�hh9�:�q]��:�������u}Y��i��0d�"�����0ïA&�*�e!��i�
��7"E3��A!���������_�Sp�^r)��r3�H�� < n�e��LL�S��������Ojl����������!&xN؋ȑ���S�c�ך��t8X��cXlxVHYEB    5e46    1530������$�d�Dg�,�?&�׸L��#����S�o^ �P`�\o��`=�e�b�C��q{+Jt���+�X�r��Hz�'��y&R�q��o��������!f;��"Kf%K�e�D�w��vD�a��.[	�yo�i8��*\{\�l��[A��a��^�D/�IzB^ԭ'U�oמ�|]1�̯,g./�L��Y$áw!���e�(�01��_�Æ������������=��ԕ�ne6-�X]�kt��=5#����t�����L��ȶ�!��c��VHT�Uq�h�� &��+'+��o�&��?KH�x8LDF.�/<��؀�7%��2�nF�Z�5/p�l�s�Vx-�b}�C�����(�YC?3}��ŀ��4��ESE��#����VL��pI�08�I�L�j�x~���ʃɒm�\�N/�i�V������Ӂ��{׊J	�bPh�l�����r�%��K����j�=����noPy?�>Սm ��<�=ڸo��4L�w�*l��ܻc1:��yU�$���9�d5�>�#��\�S��ٵ�@~��Po ά*㯬�Mwʺb�A9��Ho����V�^�:�-����+�$�1�L�����<D�Ct�xv��[n8�"$���T8�b,���(�i��I��O�/+k�,f�VG�=��dz�kF�j ��R%���EY�B����]�%���mn??�G�7�3ziE�Kx�&Ɉ�?k>�
�9E�GJ����(�{�=u��TY�����&J���k �S���K�%z[Q����3.�N�ԼwH����rj�V�]�&��n��e*��%fo]�6��/X�pú �|c�������7|��ԗYAX-����V�9Cb��,!B�>�CfՑ@���6VqJ2���fY��-=������ٹ�OH�G�Xb`��B����񜚌<�H,�ns�E�T"���SＹ�'�D4ׇ��CИ[N�����:���r�����h����T�Q��(Ϙ��	���&|9�BIx+� �^M�ݰ2aM���H�-�H�j�	�����5˿[��^Q�:�0���Tjub�#僧%^c{V!�i֫�R4���F-�ɛ,����w>6e5����_���s�~.ͪ�ǹ1 g� �,4�02@�O�a�DH���Ye��R�4����{?��L�4.Xm"���l��e9;�+%MO������[|j�zs\m~�/6^Z����Jؐށ�G sFC��������_��7����ISN���5��s.�gL\@���LI��qߧ"�q�zľ=\sŊ��]�R-�#4>a&O�D�T��\F�4W��9vޞ���CO$��߭J�4��0.5�Ȩ�;����Y$8t}��#ٝ��qFcg#7�5�xosZ��7�O(*��?I�ۘ�8�H�p=W&0��I�"���J+��s�;K�K+�{�� "Z�#g��e���z��6�������;Ԏ^�}@C�.|=R8�.!�&}a�Puf���rY��X��i~��Q&v�̐c�̇	R�-i��b��3�]S�.x���z��h[a��O����z-!c���g'�7�mmxm�J�7~�# Y���w^_6�GX
��������)�S�����1"͸U>u��#�v�.^}X;���nad87\	����BJ�a����X�?�{1p�k��/
`��a1�ݕ`̟��ǽ�fi(��^I�����8�Y��%τd�N𾰫�KQT
�?>~>Ű�l��A�t�ы?���r��.��$�4��E�ҹ���I�� ��_�%�=��=y��b�,R�� 4h`,�TSq�6�Ó%��;���wD1�:���:b��6�(1��E��$�AC0�u��̮nfN��>�0˫��֛�~¯�P��x/���̟����D3�,�8E�����s�)��r�O5I�8kգR������@6�ˢ����*Ұ@~�Y[�ۡ���h��b�������ߙV��;E)B/���~-��H�a�BO)|fi���Y��!�tք����ϕ���qeg��W�;�k�u0),����R�h1�5�`eI�q�C�9��v�I��1gB7ͥ�l�C�L�^������_����9�6��䟸��!pV7����ϔ��Z�1���i�������r�^/��p؊�����5T��V�,�D���C�?`�~F3�T��:L���ޟ�x�rv�gX4�����O���(��~oI�����:��� ��KP�le���U��ع�t�uQ��i��*�����f�����>�GD�����ft�J0k�Y/��ڽ̈�V��f���B�1|A��aEC��_�㸖v2"���]9<pwh���XsL�i��y�-tʄnc�,i�jD��B�4�?5w�F
���C@E�x�)$/�[2��qi�!n��h���1�W�@(h�G�O�m��uk���5zS�d�_1�7��zv��g�N�i`��1����sf�|���WBu�q*Y)AncW�X&�+�
�+��W�U�����t��An�?�R�;*kS���.�eH�V���ts��Fq���p�ż��x��7@��3G�(��\k��>?�:���
b&��]Aӂ8�����>3��낖��S-,�No,��z�B�!�e��o�*s%��31U�<��[Yi��d�3�,��)��u7{GW-^���\����͍�*|S�a�bU���q	�O��j��	�5�SN��ٽG ��s�<���_�]GՄSI�r��,��=�:����_�:sv�މ��֫�;e�\�02�
���2���-*6ʺ�kȎJr��-���掷<nu�S��	�i�y��νzu�x,k�J�/��0�V�&�ޖԑ?Z}5���s�j�(L�?�����}�vͳ&�%����I� �q�<>����H��7О�9�A͐���}��;u���`�?3I��xc�.�3�u�-�}c%����/��%k���9�0Dp=���7��1q�������t�G��9�U���|���R���3�7`�3B�_yф�H�b�������#|$h�o-�/�
��4�j�X����:*l3��Bq�}z��eK��=u�7M�9
�X�Ӻ/�3bvQp ����KQ��7\�@=a's /�$��v�F�X'd6�tn��5 h}�� =Ȭo,K4GɎDN_4�
���2,G��y}�BC�ah�xu�H	'�����Lϐ�jױ��I���g�h̐���	��Ѐ����k�!�&�->���v iUo�P}���HD��b���4Wj�#��s�_*�]{-G�I���x����D�&�r����X�D���B1y�^��W��RB������ٗ��XQ���p)V�^XI��( �<q?�
���5�W�A���4���:è,�qo��������`�j=��Qˍ*jͲ/�g�����/�Zᯠ<�a0!�)��a�;[��E8�ӥJcn$�>�bi�=U�����8X��X����|�4	��+f�!�q%F� m�ѦGc�/|,�1��l>�d�)���ɧ�[PK����4P��~LA3��3?��$Q���;�5!��Q�v�˹َ�3�%����Y�V���H"t����+ء�8Iu�|*@��*��f�D5p�� ��Ve�E�Rje4W���m�KJ��Ɏ����]$��($P(���obQ�5S}�1Ȓ��:(��ǳ�[t��D�w��O�A����L��3rsu�kl��^$�?�%:��l5��׆�@ŉ�Ǝ��B��$O
9����	Gp���P�>���ߔ؇NCB�{8�&E3���V�'A�A7��OƆ"OGc*Eht{]��}��5N�_�o�?���vȴʬtt��	��[�!��7�l9@���[IS�~�M&/U�I.eAC���@�c��@��῿2~ז;,���Z����^�
�9�p�G���ԝO��w2V�$�Sfg�I�Q��%ժb���C8�gR��f�FYe7%\�c������0�d�N���r�H����!Lx<_�Rv0Ѣ9��B�sʘ�r��r��[�U'ܺ���0�O,O-&+����$��4�ۧ�Z���(x��6s��U��HA�X�ɓ���P���UD��Gu	e�}���#��)��'��G��   S��y�e�l)��S��8����A��o)���O��q��ĻA
OH����D����Ӛ�0G��Q$K[6&�p�����Nuk�hA����N�f_���/��ئ��O0�.$�4�o�~�pRM�3L����Z��ʊ�X-��~�qq�1�D�)E��q}��[� ۾��k8^R������ǁT���̈v�v���֖�skY�/p/6�M�v��q�`�����c.�|�A��du�_�Z��?�8N7�P�2�8K�/QG�n%�,s3�A�灾�������<�p���1Y�J+��6R(�#_n�J��u����u�I���%�Af?��5�ϑ�4���
2�$-���L&a@Z�P��ڥ��7�^�~a4)��7}�yȟ�� �.�0��4����NJ_1͈lblo��?������~���K&��l5��%��F�9�h�D�L��KJ~%x�����op>y�	�:>@�e�C��{�H'J��i�"i)$J(ld�U����<]���>V�9p�7}�
0�G�M�C�a�(�/(��kdA���]%���>�7
�'E������~�N'�(*��h�:�9[���{=� [���S҄W۹�ن�R4���4/N���	6�i��ӌT&��&/����� >�I��}g����xR� \I�͓�~�!�珼�}7�9fiI�N,&���T��)�'К��#�8KO�08��*4>��M⠚�YJ�t"'��� ���K�X����yȰ|gvSe�'?P	���Nk��D�day^z��>�cW���:��X����.��V�*n�Y�c��Gnk��e���耷��"�Ù�?)���Ĕ���+E�w��՞�̉��3�H+����X�˩ނ��O���%a�Ii-��\�g�&#a`���KN�����h4�J��9~̘�kb<h�nǐ��ڟD��S)�S�M��K��Y��|>Nʉ]������1�Te��m>��++�E;ֶ�!�qj�(��P2P�O����y� �;�X?!3Jz�����BF���tTuI	�(|�_(D�-��K�W�:s������1���*�w���8]k��5����g��Ҩ7����k�^y7��`�#)����%?&������LHMr��Z���ُB���]g�Tp�Ⱡ�F�)�X�����!5�ܳ�Ok4�3F�9U(