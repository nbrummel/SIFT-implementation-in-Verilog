XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��wDط�9�I���]W7�.(�ʥ%�D._B�l�)�Y�N�,R��_�,�`�	�wr�;�9�.��pv�����0�/�[Wl��*.�P�=xKT��Ӵ�����!ov��D�@6>�8����%�Pv�j��k��oϏs���ij�g&����8:�(�>�R�>��9z����F�B WC7��u^������$J���#�����+��G����k�[ v�g��d��\:��0���^i��sV"0c�}��E�B4
�Ax�*�J6@������o�4&�'>?(�	�H�0��.6t���^�$n�>X0_0 �!���Ǥ���")�\���
YZp��\&'e�롦�0z���p��u�'.~�͌C�s����nj̀wg�O=χb�e�2���}�̭�u�R�>����� ��� d�,�m�C�FI��\�QEhf@�q����ód���fi���d�g�p2�,��dZe#6�ةG��<6�q�h�[�wJᣋ�!��c���e�W�{W��0��N� +Bp��n˰��G�r�j"� �9�K�h��\%,u��KN�f������B��3y��\s�ĩ\�4��:e7��������hk���d^�֮xJ���Y�>.|�e$�{Ӑ��<���;\#V���(�l��GWl1��}3���b8_Ѻ����j��gW�Gl�\'>E�.�eڔ��Z��Y�r,V$��D��VڊQ�B�����1�H����>cq��@9ђ��XlxVHYEB    2fbb     b70��jD��M��b=�j0��9�^��k���ͪ�����n�U���&�'�Y�[���3f��+�ݸ�1��?�(I��Z��=a�ָ�K=?��*���?�fѾ�vG��Pk�.��d=��/�zkJ���)���y:�:��#�N�J��D��
̊�æ����<_���m�s E� K�Ʒh�6f��;�n�^��tq����kH����]�$�_�Q�Ѳ�������U��@�c���~�W_!W�7eG��"������膴0YbAqj5ed�nH�hkF8K™��ݷ0�Q��k��P@�����Ixx��%�k�\j���;�v�ۀa篃@��&� ;��s���}_���,����NN�w��
�a�l��˄؅�iSQ�P�m,J=�1��#�Tz�X{k���w���o h�@$u�Lh�ѕ
�gF�g9a��Ǝ�1��\�l�?<>:1SWE�'�������SۂX�(bA-��|�]�>Nݜey:6�^T��

�����}��4���H]O��+�-4?-n��y��gƣ�)gL�.ӔSى�\Z�a�vv�K�˜|���4%��Uh
|���?��2�Ёߩ��a�� vS�foV!��h��ʬ���Xzk�(,$�$+�rL��0��o��W�X��>����+5~գÿ�_5��#���^� �M��^�)�$��z���w-�	/��-V?�^	�m<b�bS�b ��)2o�ǜ�,q�r���/8�D3��7��>%�|��+Qa�J$��QF��A��ՕD�t������֬S0���lY~����1��@��+�C���2Ѣ��"D-$~/�[�h��L�@K2�z3L��
�ԙ�-fωQ>)�Nz��7�<���/_�f*l�`O�����a(53��dI��-�Y��wG<ƵŬƅ֯ľ�R¬%<��F9!��b
�Wҙ�vY�
�m���H6��{y#SќVΖ�0@c�HKS�o����~8�>l��	;]P[�\�O$�Px�Σ�ՙ��3ZKgN0Ѹd�b�8���1��������,?��]�T����fN���&��$:�i��C�o�2����(M>?��f���p"c�g����A-�.+RCo�ko"|{�����F.���- ������
�c�kՠ�-�[3���z؞':��E�lO<~ZA���-��2���4ǭ���G/�,-s�Y�dc�Jڜ�c�o��	;�>j�x�֒��^��Q���0|�������]�E_%�Ć�������#5�c�%�^/̝���b�%�(�i7��!�Sde��4��M��T5��"<�;�}>H
�G!���-�<Q^��f��Уe����.���o������׷�_F"��g��Ms�����co�t˜^��LN症�W ����͍��%�@	�N�3ySl3�2A$Uf�䭭�����E�Kc�Vגk�i3J`xg$��>v��=j:4��)��ҋ!��	M!����`�.�V�AʧU�M�?@�,
��E��j����G{��ƿ���j�#+�g�6!�5=���Z�X�����5<�q/�)����vG/�>����R�?��f������<��A��l�JP�RؑER�]?g�l��	ߵ��&d9�J�Ka�-��4��u��._@��͢އ�P>�N�2���u.\jb�%x����Q)uoA�A��@f�'W�a��P�I`�>�O�J6�(�O�<x���v�0��R��.�2d�-�����Wg	�c�k;����8�PA�/B����j�~�'�ht�3@��?��w荙W])B�P��ꑍ&�xי姧�R:�o�Uh	���1d��w�>n�E1-h`�wq�	�l�@��D���`�/k�Σo�g��l�h�� #��V|�)�=S�����LY\���`�j�e��DX�j�P�[�$����M��
��5P;~{��1-D�{m`�ڭ�z>�$a�k���?1�>�8�$MWy�KH��@;���yQ4���8��V�&���M�;��#E��p�n�	�
B���Ӹ�A��Y�7N�u��ga2縞c����6;�����Ԩ����'֭�YV�4x���jsF!+�`�;$�D���������Z�9%�3��C��k���xB9�?7D3�����.*�g��c�yO��DҮǇ��B������ ��4�ҧ�V('aN�ZH���D�a4��^W���$G���`+�ǜ��������G"��q�	eb����I�l�s���$��
�)�cc��82��$L�>WOB����Y��b䠫d�_����l="�
��,�?��3�d-4�b�>�ۻ�_oi�<�r0�e{��i� 3��n�9�D$ލ%�gέ����o?J6"0;(���D=����DP�"������X]��s�V���F����X�Dn��gVͫŉs�ު;8�"yt �7�v���jZZ('(��F�exx�Xb��?�]��a�S$��v<BD�0m1��|`	���6 ��d��Ǘ�TcLb�$�p�+�3�P Pd:�%���	@�_M�E��g��D�"��%�vpu���;�b4r���C���75� ]��(5��l}�&� �G
�����U���.�o?������t\<7%0ϼ�ϞO���-��x?��^�(`u(ĺ�=z٣Q;�0���:���[;�|��� �ُAr�{���3g�[r�L�|���\���]F�R���`;/���,����h�;�7�5����V����1��6��>
�˿ΦS�h6�`�͝�fU��嗨XI8�Wi&8�V'+�A�&}�MN6��ܸ,�%"w�;���&�)���[)-�ɒ��#����.�N��7K-���a�CG���묷��4�UY���J+�����;