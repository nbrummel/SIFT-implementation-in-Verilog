XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x���Jk���toY�y1B����7���l+�r���x�~:�F,l�J�Oގ��3�n�9'F#,��jV�����(ު]�V����_�w�T��O�Ne��`L?t��R��x�a3�7#2��l��Tc���'~�滕P*�Q��p�Ѝ��I�Os�HՉ�<�����cA>C@h���A��G<N�:R'އ��h�V�ݲv��L�z��_Ai�������`Y&<���f�6�R�L"�*7"�q��u�?B�^��\�1`��H�,v�V*[�$e�Cf��J�+�F��Ϋz{��>e�k(C�`>�x6�,�X����}�	�j��;E�ų�,z"A;�P +t`�c���9���?8�ޅ������wk�j�	�Ӏ`�j~��_�+�^�gT.�Ʈ������/�sRL�D��,�b_޹�en:IΗ� �0�6���	��_��8JGt3�%	-�Iy�����>�̡*:�cP�����o%�_����#��V������17�j�RG�ǒ4?2���	˅���֊CCU`��(k�7�����AƘ4���.�9c�e$�C46���:��h��9�D�'3:�Y��-�`�1�dT;�� ¼��}>L�9�4(F��+���~tdd�K�Q���Þ�z��|w�Ç�WcV�|��FRnuR���J
�t���RD5 �1 ۸�庼p���Y������'�n�8��(<��7CP�h0�sew�r@��6=���e,��x>�U�d�v�ޣHXlxVHYEB    fa00    2470�Z��}�y��F����^LH�	�aH'��\�OQ7/習ն�]mge��G��F�i����FwFp��}Lq��Z��#��G�&2� �S�i)$���IF2�d�����u.\�q���3��a�ȝ���l�8sO�DJ�n�_�/ ��_|&��%)�$>橥�v�47O_	Д�'�so�A���J���vF�� z��K>q�M�еi0���b/���x^ğ,�[EE�� E0����f��a/�O�p��g��q�$��%挊�S�1�G��|5%�ۀD��;eyN]|�Fݏ�S���n�	�����`ߺN��V�
߄���u��F|9�{�!���N�PB����b$�P�`�x����TX�U#C�b*�iU��'��GϿ�14�x�hQ-GQ5#C4-j��֗-�7�0	 :���𜀇�{�3R7�RM�~t�F���� Z�[tBw�(C�����g�^&3��u�Z�Z&kAd�+zʙ��ڠw7UAc2"�?�R�F�d���/���x�S�6�5oR��L�PO�]� ���%��|А`N���;����g˖/�`�� :����ZC�Vǁ��C��Ds �=ӬL�t!K��fVq�η]�~$��`iF�?a�b<�YF��pX���S������-	1|���Wu�����G����ɧ����ϟ��ac���9^w1�6�)���8?9$��Fn\hޖ�A0�>���I�&=Bk���(c��v
two�>Մ�������9J���*U	9b,6��Wp</�H�0���J��i��1s�2�ЂL�6�)X�[+Q,��E����s�����y~m�~uT�['N��)SZq�8�hj_�P�g�c�i~&�c���"^���e@���rD�TϺ�jA��0����є/}sɨS!t޲g,�
����Ŷ���F>T������	��tKY
⤈�������F&�8P�d��- �r?��S)��g�0rK��n�\�IxP���p�F�O�<a�p�ܢ9I:6�|�}˻�Mj5�+�I�rpj͈vd�k�򦤡$"#a�'�d4�qp��h�оw�r°{r?)����m����iz��O�qm�w�z������'���ߣN��;�>Q��v���)�^�\�eƷ��}'��Gw��}�����/8�Nk6�_ �oQ�ӤځN��c�:�u	��63w��{���D�_ss/7 {�n��VfZ
�������M��Y� �,���}�7��G�ɸ`�
l�@3r�t�e�b��wU�ߜ�Bƀ�@q�.8�Z�ɼ�F^"-��3�ok�S(`��RSI�}=�g�g'`�tk��z�UU�k� ?+Z���{￧��@����9�{W�w�b�����q�w����F��e�7y�I�Ђ��������"=h�R�����M��~9a�CEE���e��r?��Q��ʉ��?�܎�3�t�����j{���Rǁ����ҍ��k� �a��&���ec�(\�/(V~Ȧ.w_��=#�]�u4~^&T�O�r���,G\ސN�7?9��#n�Q�5=��-1D�w�6�;�0�/�m�����o�Dk��N[[�E�=��ʕn�I8a��˂�4�&���)۰Ȟu����ؔ�(<�R���Y꽇[��c�}���n����r�i��&�	��0�e�-�C�1t�P".����/�XK�+� �N�s\1\4��?s�6�$�@-��$��Q����p�%����ֶ����A��}hT5��"ԩ"҄�b���ܤu�ڡJ���Sl��X`/���e�q�{�e�ʯ+ě������-�����陸����e _neȬ���'�Ɣ�{��<��7]��e!���S1�of7���M����[qW4�p����8,�Ұ3����ߏ����ٻ%��n�=�>�'uN�Z<oBف� �ɐuuC
FH��ѿ��q�\��������-5p�I6?|�+*|�j{�A�Ė�H�	��Ǚ���2�?���GMsC_�������1��Z��9J10�3^�
���>Y�G�LBۮ��r�#{`2�F-��Ϣw��M�v)��c��_=k=y��Eq�F�"�_9O�d�Sv�'Wz'W��޹L��mm��|����q�����t9j��3����\܀}�zk��*tS?G�,PT�_B��_���B`�8?�닌����\� DɞO��@車)���xe�=7	����+�n(�/��*�̶��:o��0�Ͱ���'��VVoZ���T�e
?AL~����_O��l�|T�[��.�ĂW��& hE�mC�6E&Y�%I[�~��*6:�F�x�C��ߨ��a ��`2���DC�f������t*}����K wП&�P~��lvn�qN6v���Ǻ�Qe�G$	�|x�k��ۮ��_?�W�H{��=����G�K�PL:DU&�I��X�'7?�6�j��ꋐ�(��c�K&�YP��>w-(�[��ڣ�,wtd�Dˀ�ِ_����C���RԮ:��P�$	�e���q��� �&����	FbA�s�,{@*���C��>��*�J�O1������w0�	������L@�� ��h�gw#��xnx���A	����2Ä5�S�̃�J���y�u�~��)ǋ��z���M�:������zԻ*�ݏ���Pv҆��*-�>ڹ���en[fc�Hl�H(ԉ�ݽF���z��Չ�S�������Tʴ��qzDVv�Vio�U�Ʃ����N�y>����X+ى{���\���`nX/dօ��z���#�Z��S�\��Jw���I�d�y�y�(�/z��� �.��L��R�('/UXg��kH�ps���`<1��bG�p:�����)�=,��9Ĉ���̕Y�֡p,���zM��:�n��`�a&��s��W�M؍O��D&�]gl�+z3	|&궋��ɘs���I�f���;VÙY|Ue ����g����[��ڞ�H�,�q�mˣu����9��p�1V����B�2���D��* �Nsˊ������b�Y$���C v$�iBIz�"��O����3�ѮW�G�X �{�>)�,��nWo�W�ca�+���i��!��������]E< ��G�m�dn�eP�����B�0d6�PX��dl���!)�7��L�k؆1���.Q��a��T~m�!ǩ����WD���ec�`�'`qa�4�lvA*���qr���H��].�D�|L�F��<z-�� �XE\��<�~�\"].hQ�s�чV�~>�7�/�a�	<������PV|���Ni@C2W� �47��v�Uݫn��N����:ɍM�@ӗoL�Sz��n�j�������jH��#)�z���>���86���y���Rdp\f�b����'�tf�*is�#�޷
�.GU��1(F�9�)Ij�uc�ޡWIH'Qc��5�v1&�K�w��һ0�b/"���.,��/��R���L8(�ɝoQ��9i�eG��O�{�Vy|)Z[~�/X�
��O��l���������(5BKb$�EB7;����:[�;��\�o�]/����{ZS9	X�@�^ejC���v�m ��(�/�'�2b�љqĸf�(L[drQ�,���_��������ad�a�Hф6�C��7���p�E=~����񓲮�<�=������ϺCu�wI��b�Kޘ�Y9�`�KwA� <���o��|���B\<�H�`p�v�(-��Q�LEF���X�G�]��!4V�0|�]�uϟb!J[I�Q}>g;�f�xG�$��a�r�t�EѿS��xUN{#������F��^s�>ѱ��U��Ⱥ$P�zb�)��A<5{Pj�R^��&���yu�o�/��+���1����\�����R?��!�ߓ����I��JW��!�	��&0�<U�O��{��E�p��L�j��,߁�f~QD�H��ߥ�:��L�P�D#���ޓ�ƍ��-������XNf��L�Sh��H��Δun�eAY)e����3e�|5��v��u��T,P������|��:e�&cq�>F�] *E"��-M�IA���ި%����w�Z�ӻP�.j��=۠ѫP��(޾��tew�'.��!�k��m�5B��?�t��@s֊Km}�{T�����r�e�9�����!,�%�{�d&�"~v33�?�cY��7��rH2��S(��	��>ͪ/���Jd�m�(��:i�<,`�T�k�Xc,�PJ3 ��/Եi	��K��Nm�A�߁�������L/��?f'��?�u����@���`Mۃ���ֱUǑ���l���W�v�Y<�JK��@P��)�:�!":����I�䘶|�	!5��#X,($�f���rٍj
�q�@��'/�0�s*��O0��u�z���*Y2����uQ��{���M�K��_���f��%k�l3��ԥ��k��C�%�U�W ط�ZU����(���A��V��U�L,ac��]	�<��V��WTT�Q�7r��#a�#������g���VXk�8�ܵs.T���[��! 
>}+0zo$H
k�nEsۨ�b	 no�ӍӠmQ�����z�E0e�S� ��c>�
l������^��SFv9ƒ���ڋ���Qj� ���<(2}@�睉�yWNf�}ɨ
u�Ǝ~[L�G����bG���T���l�h��^&s�RhP��(�;����j��X��j>�]�Eq�����Vq`-k�h��+�yZL��ťk��"�~�Y�`�H�`Fl+�!gY���\�X���%%�g&|9�]*i�t��.�-��PŰ������Z+�x�42�~���ܽ����{���j�kM�u��I�,�w[Z�2ym�h)�{ tV���U����5���n��d,�a���@P��"u'�ځ>��Qѭ���	�G�EY�����^��?'����3K7T�n38��/Ϩ{��b����?�ﲛ0��9<em�� �8w
Fթ?KO#=����D�ō؝���H?X;ۓ��r�aEOlu��Zє\:�G��iQ#�� t2���W6�b\�)�?Lzǘ[�Fww�����;!6��3ɐE���x�*�}����H�
	��۴^l���8n��0�Oޒe���'Ȉ�-�A����̟���nݍ��_,�Sttf�ً�8N��9R��@��FW"�x�Z����X��"�;Λ_�O'�f�xT��A*��
�|�d�����n���������y�f�Y�bm��{��b�9��B���J���oh�=ܖ��/�K&Υ�:�2��3V������H.aS�\(��e�W���oWj���rT�[kq�+N�kr���*$hS�q�y�Z-��C���Ր��F���}�׈�,�:>8"�@1F�oɉ[��̎��-��E��/��9���ęS�0M;eo�����y��өV)��3KR��P��l�ӕ��b�&s>mN"�Q��&"�D���!n�s@ �����c6ݦ?$W)�7���~��BX���4�T�k߬��x�jB�?nhLN�]��CJV�SdOt+��~�*G�3y1E�4�G.9���	�R�uQ ��������l*Ǹ`�nO�1�.Xi�7��On�����T�L�-�B�eڜ2�/��<��k [���4=i����1{؆��RT9�E�tp���q7K-���G��șT�ue@�t��v�^?Y�b^?��/H]�#]v9r���d��Km�m�(�GL_FKiaq1���蹲��<U�64U��bπm*cmuj-E����L�#��+�%^P#K���E��H��h�/�n� �l�չ���6����d���R�Ui�O�����\���5 �h�'���6-W@�?�� j��� >�9lT(�k>yچ`j%}�"\�$Kr�k���@���r we���W��D\�qi ���?Z+��<�T��w��7���5*��h2n�eIS@�dU`����:�mL��02%J��ǰJ�Pԉ�o��H=���m������q:(b��#
>���uQ��CMW�]�>�~-��C�a<�B"�EK�ĿE	�'rB�ud�KFļ��뾑�~z}m=7A�~�%�nm����#T�����\����N�Τ�t�u®G�5hxi�p���<hM�3�^��.G9C�ɘ?��@�0ޮ:�-L�/^Z8�T�퇠t��Ei9Rv�q������T���)@G1ζ��F��-����Cw��C|op�:�AL�wv.���sf`�yI%�|�sT:bI)ҥ��ta1����I�u:�x�L1f�[�I'�Ŋ�P?�N�O�ݳGV�1�H��ϩ{K�
@~��M"��}�`m'=�������}M�yL�Ǡ	8,d�m��u�)�[�X��.Dul���A�@ײ���Ƽ<�;*B�Sx�݌��Y 5�}�酪 �g_EVe/��r�pN8ҏ�EL�%h�D���U�F�ܦ�fި8��e�d΂�����`Ks�6*�G&3l5�ڀHސ���峵}]C�s���upCϹ��V)ʈ̷'s�L��v����ɚ��.}\ūa%���ޜ��qe+�p���ӕ�8y�zԮl1��G�#Ǻ�xA�j��{�[ș�v+����BP�ߒ:ɼ��|-+�	M{-�|ˉkS�1h���z�u�g'�u�譌��4MJ��>wM���Y.�̵N�i�#
�/�AZܼA�u(s[�:�ڮ�񓨃O����i�{$`ߧ/6g�1T������Au�4Tn�`��W���N��]��X�n���wܺ6
��y��e���ϥWYm����6��=����Њ�Cse������+�c������vu;�*X]�p�$�}�H����=��`\��mo��=����]�����L��=X�������
BV�2�{Q�`�G&�ԫ�)t��̦JP�^�Ko2}��b�~	a>��X�|������1U���&q�n��� ;���w/�]���>(��$_��UAh��Ay�������8F�-�)��$B�=X:~k����Ŗ��9AD����#ÊX����/_�EhJ��,�f����YiBw*�+��Z�!�W��m[Zx ��1Zr�eyeL�m4���Z�m� ��� �+��na���|����������e�-1�����ި��<�'��1��0YZ�]�C��k�r���"���6��t��C��b�lE���<NCJ;��4���wޟI��:#d�ϖaA��X��������	r
�}Ӕ�q��E�z�ʉ�$�!@��0�A��/��^.ʬ����e�1��=��?�Ɋ�����o�
 ��c[M��?�Ԅl�w�0à������5���%@���u���޷�D�fG:��2�bil�~pu()�3���7}�XN�� 6ѭ�Ià�}h$K�Jp�y¡�(/i���!?�*aX�!��W��C����h�l�3`@�T��{p������Y�h�T���u�o��N�d'��@�ؚ�@k,% ��тq`����cu8f����YG�a<��Y��($L�Ks��azԊm 5,@�UPt�C��1��ֳ:OV��@�K����YjAeQE�i����P���?W#�#��Q��oڐ����oo`��.�� N�&r�hX~+,[��`��m���55�o�2����}z�k����)z���PjOHJt,�,�����^D���ۼ�Gjq~����M���#�7���b_$#_��,�Hن�(��[b0<�SJlX �ƴf��ֻ�7�8���|��ZQ(�]��Fl��K׉l�di,�Н�A�@<>��g�.�(r��#Ƴ���f�h]k����nA&��wēq{"d����a�����q��z���M�k�1��#��Uv���+"E|	�"���Q·��K��{�G�ĤΑ�V@� �!��V-�h��3��`���c����Im��.G]���K��,��I�֟`��جM�����:%Z��|]E��X�a'c̷�ՌE!�眞�FQ_�1Q�Gk� ��_,��X��Qz��nc��.�g�wxj;�����!�#7O!��Re�:��H% �m�i� l	��pxs��Wo/@���ZX�L�I��^��6k&�O�S�Qp�[@�{1�QޑN5��ٱ�I�z�����!��9������
��,�FmSx) �L��6)�#���St�)Ԭ���1��r��I!+����?R1j\	�[�Mb�#��݊JX~7"l	٫y��x�Җf}S=�-ދA��v�����ޭk&�/�G���aQDcai�	�����a�#�Ԛ��7�&^�d�֌EUv�^0�!\x���K�	Y! �x�J�  _xtO,�6S�����`�m���)r.���Rd�T�''������|N����Ϲ�v��h'}	�POќg�����繓 �)|z2��(���荪X
�6�:��~��p׺�d�c��y���D�gML3SΘ��5����®q=rI�LR���a:�osq6+VˠR[h7�6m�<�)ݬ\���Eh�����\�\����4�i�N��*���*�^�I�Z?HcA�O�ȃr�j�+�G�����ck��������ki��M�FYT�E��7���_>ݩՖK{iF�/�0C��c]��h���`�u��TcX���4��o�����[?����ץ�����0�8�ߚ7d\PH�.u��eJ�(�F=�M��Y��q�C��vV�K�u��6?�i7��3�+UϿu�	A��o�+�'DL�r9����%��`�rg��1mG�hX1ɥ�����D�[
Լk�
��0x_u��XY�������%�	����ÎN�g���ް����4�vZh%;s�ǘ��]N��9z���E&���_.�;ƿ�����͞h�*��`φ��O"���"j<��
w���L���?��T�Z��H��y"D�k�p����N���p�N��'��gPB?"��o�|O���X�"��#+�l�K�v��)Ȓ�d1��c�{�IbYOFU/@��E��/�4f��A�w��2���0d�J�өK�@� 7�����d&H�R3�	�L���rb6w�.��=|Ð�4y%L������O�BM����F�XlxVHYEB    fa00    1b30ʣC\M����̦.�?�x�K\�[��I�J�U-��
(����i�5ϩ4>uGh�9���!C�g��{�r��*J_��VZ��vZ�x���E�$NJᵲ�R.�]���K��e�'�#0!g�AA��Ǹ�������,�_���8��kRo���'�^��̭Ez��{�뱸��Ԧ����i#V����`r�U�q��m��p�����+Җ�2��
н�C�G�H)�Y�H�}SGUN�������c�H_�(e��NK��������Qg����;���CV;�ٿ�tJ�mB/�$���|��
0a���I�>|�P��W5x����Js�ghM�L�xP�t���+i�N7r���������)��?���)q7{,R��;ݺo[I�&�W6.n?l���������G,S��ob�އ�j
gCl��j�PV̂vNm9Х	��:�򟉭Vț���8}�ݡ*[�ɤH����J1	��1���]�`,�:"`1[ �j�:<��3M�ӆ��PA)=3����r��g�M�Y{d�vvseG��?�/�3��~~(-��C�I8����,��� v�6&��;��f�"O��s��!�uc���#�yz���jx���P£I^�4j_����D�Z�ֶVaw��ί���<-e�\�&;GRsP2}L�����a"�U L�q�1-��+�PhM�/�~v�=57 o�l4_q�W@]�<��"��9��`f"�+R�X%W��e}ŭs_ߙ�;_|Lv1Ý�����%p�Z9�cU�r��^Uy�	�6}U���8�OU�o���o2�N�A!�_��]��J��X���W�n9T�R2̉��	x�Ϫ�G�&×E%U�����ی�m�k�wQ������"��l���bMw�����L+1HTV��  ����s��ZB��/%��Q$�S�k��	YL�0	�SB.�Cy�+�y&�:����Ҟ�%?�:�n���P���������(r:����q��%6"Ja�&��%w�4��fht���5[�(�5���0��r N�F��rP�J1"ڏ|���~��Y~�t-P�O�4d�ԅg��M�3r4v;;�0��|�\�����NuI�f�����Cp�,<?�:T�����-����_��Ɔ�jٌRiŎ�1@$?qR���KƂqN_-ЮB,PZ_#�-Ŗ$�r�ޞ�����d�Պ�?����8�n������N��5��K���P1���C�+CyJ	b_�-*���}�nB��&T�ꖰ��1A5�(����!H���&�	�q窊F�?�!`*2o؈���#C8zmKL�6��M��!�# �>wз*�+�NN$��͒|�����q��<��!p��+%�~�	�U�R��D�%�c�vw�.p�d�'d؇���.8������<�O�y�ĪW{0.�g�8�"��GViEy��~ �!SW	-�v�
g(��t�of�4���n�Z9²�D��>åD��C���E�-���vH�
y6��&���O��2�m���9�Դ�t8b �����mw�������_��=W�W����9� 9�8$3�$kphE@Jǫ�,�a�.^�wj?��C�dà����˟G'f��`�섦 �Vw\��4b�)���[�\x��,d�tX�S��!T���$�J�1�ul�l���z�z���2q�����c�����PO��m�:�D�}����i�J����P٠���! Pv�`�e^�}�B\Ŗc�Ԫ˓$��H)�D�j4�����Q��3 �Q���H��_���9�{�L.�-�5G�ם�)�SgV*-�EB4�����1�u��R\��S`gA������fH��ЖЭ�� =�� $х[ �:"�NM�s��4�γ��Y�,$��-����&@�ZH�'�1w:aH�j�u�+I
cd�Z��n4�e|�A!`�o��'t��G�\6XC�C����t����)����ލ�&T�l�La�<��}�hU��䫻]����l�r�u���a��ؓ����v�Q�Z�uv��M���U��js��I���� �u�6Es��-�7����T��j����h�%S"��f�\0�M�י���4^7Ǳ���V��;͑N)vUX�q/��0i�����%�������=�	��������	��_q�m�U��I�Ռ<[�s���$:~���v�շP�%�e�%�6�&"C��,\kQ��#����C�����t9A,9��U+�L0��lx�Q1- ��M8��+"a���4��r�3���&��Y�5}�c��?��죏He��3�s�m��'���<J��T���7��`�ԩ4�x��|'���iV#�K1W��%�������P5��T�Ȟ���/hiy�K��e%o� N}@�~ym�Z~W-GW"�]?E��ɖ
p5����"b��K}fx�d�5|�������A�2���5�O˝d`�,Nzq ���ɉd�1]y�l?P7�L��w���Ȃ�8dgތLΗ�)G�1����j�C�^���M�c����'�c�a4 
w�D�$�N��3���(�@%*f	SJk�����Cni����]e2{��S�@�M�f���Uu�̟S��U���Y٨]��@���Q�Z��!��I`�����ڻ�O��aΉp�5
8*.u�h=��ZĜ�Ȏ������=���J#޴''6�Sl&�fJFI��D��;8�_1~*��	u�
�����I\G*>
�m�88c�����i�5�'�?�X��H�\!Np{�!>�����c]/�$�!$Sm@�z��N��g	4���r���ʛ׉�"�~�%۬P2x7%=-w�y��
l��t�}�
N�U����7�L�#�����T�EFH]��)�)���z3�l��zbi�.�9���e��#s⼳����G�=�5�����%
2	쒔�[���i� �=z��ZѨ |97a� t������-�f%[.�XV���c��h-4_��u���+�����?1���S�)a�gc\��V�:��{���+Q������D
���@����n"Y��N��bLh��Ac�O���zgk�-��"��,���T���M�!�	�����!'��"��Ju���Ʈ�nD�>�x��0�\��_��E�ȴ�����
�
����&Bb���5!.TZ�uH�=�cw�&ѧ�ݫ�/������*�Ʈe ;���Vx��O��� |��mx<pZP~�cFL���e�4�7Ib�!8}-Q��:���&��IOX�ŪI���xL؎�l��Y[nN��q_N�Q@ ʬwᲆ��M��ԄBE�w/��i�������ު�2��D} g7���T��р�'�eR�ȣ�pm<�<$��޲�	��?��X��Ln�8xc���Z$�6
C��t�eIm茙"x��u�4����[�m�Z�x���ܗD�X�I�9�'����}ٴ!�?
Pt�c����9>N�Ɏ�<��ޭ�1�]F�;ֺ���|+��FO%�լ������>Db�� ���O��S&1B�j�F�Y�i��(.OI3�%'�0�������i,�&@z�����z��w1u�$;R�虵�
�kl]���,��P�5��m�Yq!4�T�y	]3�4����M������O�_e-���aD{�ZC=�t�񳅞���}�im�]�4HnA�����Q-zsqx:��)dH�5�ٖ�@��Az�N��a,�a.���>n(�'�1��8(�o�	�z��ŭ�E�زB%s�Z��r?�y����N\�i�
c�������l8�j ��ש��bh��6�?��P�a��ͰJST�e�*&	��}Y�9ZY��R��Ş���O�]'�%��\8EE2e~���ɢUJ��U��n�ꃩ���P�f�څ��B�ӌ> 5�I&��(�3^]1^�_�N�`(�p��k]�M�e��u��8a,<}��Ρ��)��P�-ߑ��kLC!�ʋ��Βg
����D�Į>ca��s^�6��mz� u��?4W�'j��pG6�ŘG�S��p�3^vd�%��q����S���K��U��Q	�C�n��|���>�������/3����`TLg##��nP��h��$y�%n~�f�n�W{��_�	M�(�Q�t=�������Ä�1d�\߉�8kyh��h27�h���|fD� �I(��t&��YU�s�~t�,_�����[�B
���l�J��J��3T�`!1ab�V'shqKJ�R����a�GT��3����������x_�����v}�ڃI&Ek�KdM�F�xk�2K� <��.r�}����O�ezl@��y,Wn�>QS-b��a�].g	�� �ibk
yp6����e($�֞��riӞR�DKJ�#�C�k���dv-�U{&�p�6Ŏ'8�v"z#���1��?�}@6\�/G=��9�-�%�l�Q�[�����~kŝ��`�#!�>>�k�e��N%𨇨�Y���4�:a	�ӎw���tߍ3䔅.
e2=�ܗ'�`;�԰f&J���lÔH'۬��XH�h���o�.�6Ϝ&ܬX>���hg Gh^������)|.�_�g�Y��R�B�I�}����U�Y���w�C��J��FK_�im׷#���Ku���#�L�K��|��m�*!Q���oS�k�"(�>����L�HԞ���ɫ�U��w1�a�K�J���P�e8wM���'=��,��5-��F�W�3���c�g��?��@��5Տ��F%��Z9�z�8��P��\�65�����Dٗm�s.8Hw���Qr�J��HV�s�����J -�d#*6XxoBα����[�9�d�5:N�_��϶��ma���?3D����� `��,�.6]�y1�0�ݒz���lN�|��n�>�E����b��ց"��3��q�����&|�ѾT3���b`]��Z�:�c�j D�4��}��\��XXq�nv�4d�P�e]�I5�v���B�mZ��?����_�y�)�ۃ��X5��I[���?��\A�s&�ɜ�^i۫2����*���޵FSDZ�KEB����$(��-TZנC�Ĝ;�4P�D�\e��ɲ/��Q��!��wa.� ���c���:���I������P�-�ͧ8Q��拰�ƫ�\:'�Xɜ8K%�7��0o������h��w�u�?����?�J(�����vղSέ�c8����6�VUl'�S�NE��TH*sg�i�9O�ߠ�L9*]e���D�2���v�C}�xmn��5�wc�b��Ԝ�r�H��[:�ȬmA�%�Vƫ�F����˥�?����<�όҺv��:�p�jP�{���3%���w�q:N?����"Q��΅�>U��\�K�f�'ZTY��@�Q*m��>�W�o�j,`��YA�p���~�fI���<�ջ���o�(����m���'�s.*jVc,s�F21�a��;<:Uҽ�~9*�:���|�M�M�R���Y�>��'+4PT7��t�`��(�'SA�ߏ��^��a&LO{���ո
n�� ~�' �P�W�UH�T�ү�
:���}$�sE�ue��!y*���[�ɺ���^g���we��o�U�?o��7?܊�2�~<|ʫN����]�<F��R�{[=����M�Zأ�S�2d��k�d��S��ݲ��i���S�Sh�����\�àg��2Ѩ$����	C3��xM/[�oRYb��>���J�Y}7�i�D��H8n����<�+��,�!���\p�i$j���kѬ�'�x �]�>�n7̈��r^�)o.�&�<~����i�|��7��P��/�!��L4�*�&�s��H��I�P�W���YxE3$6򣢻c�y�X�B�g�i &j �z�nv��4?��n��ʻB�j	�ep�|C����c}��<����a�-�꼅�{w�����@p#W~� MRXv�D1w+�� )O?_�g����(�4s	���}��48�DC�o�RuWP�1� <���	t�KL����Hd�3����{�ܝ�;¾�xL�u�7w�u{����T� %Ae]��7�Or^�L�:Ɣ�����-Ů2�d�&\!�	�	�6K���#�����ze�=��*�:��W|(�R�2�r%}�)b�E�-�u �=�v��(��%�%\�X;�3D�-]���������Xl5�nQ����2"W)xY�cBu�҅�މ����[�����,�^c�NA�^�g����+�P�u)�W��0���H�[�x%�|��{D�2�L�`����Q�3�,�����זvd(����c��!C%���F���		���U�	��S0ٕ������L�V/��Qβ�~ `��^���pyo����>�P���C*�&3JA��m�A�&��/mv�2�����e���s�3�Nս0��K�I�ua/���|��iR�������(�!Igb�K6>�A�-lBb��CZt��"�������J�l"�Lt�;ח⺌�*e�*��J�6%�b�omGlCH*}��3�y'5����ng�3Y ��"&��+�[��s,e����ܡ��P�
S)���v��m��k�U�Ut�R��6��,<�+{���%��~�����<L!�)\��5%ɘ�'j��TC��U80J`F��v���|��!�n�H �M ��x���<:�@G�������C���NCh��"X���|8n�N��~���u�e�91�ھ����CL7Z0��6�ȏ
��fJ�9�Ӵ ��*�֧X��AA����k�%��w��d��w�@�#��a�w���XlxVHYEB    fa00    1950�ã�]faBgt�c���=.�43e��~��3�T�d�:Đ�f���=�ٶK��;�8�����C��;u�{lM^�;U�&WIc�M�aoW�x�>�At�-'�)��������z�n���� >�D\�[�ȅ�6Pz��{��3��%��A�<�BGuC�n?��Q���$�����0A��M���#�M��!�~��a��Oñ��TT�}؊�>����iF �*Y�ӿ钆���Pi�U�e^#��p��� �0��~���qX�e�&k��{��O+(!�N��WH��g��0+��"��`;r�dy���^�P"���^�M	����&�[��|Р�uD����
~��F�#S8h���͝���a�9�(�!ge7zs��n2��v�	7�?���^�_�|{;��5]ǕD������!_�����v���u��\�G�G�P �����Nj����!���""��ex�����\-�.��n��H ��1�4w{0yX��EQ�X�ܟ����QH��] F�6m�5��I���O�r�F2qE�Oglѳ�XhG]g����9u�=l���0���5���BRS�.8>q���p�m�Ҿ��4��^��p�2ŭ9�
k�i���7�b��T���b�L[���<Yy�}������~���V *�s0�n
{�U���s�O�2<N �&�;Ɵ6y���;f�j��o��p}���\ȆM�8$�l5�����R�%����b��I䛥J�P~ջ�%y!6�3��'t8��y[��x�d#-j�-�^���.#LN�D # )4�����(�bb�[J��8��t�Pк?��j,�$vW�^hDKz���@�>{�N�b��>�%ᇋ�������� W�E;}#��R^����+�.�,Rv��~[��]���z1��x����#`۹xȱ�:��}ǀ&� �㯸e����U�iEÖ����OZێg�,���W��D�U�r�p�S���e�y8�c�H&K�;VF�^!�#-[�׆+^���bP�9��V�l�A�陗D�B���Q� \�e"����X�ѵ�I��DX���u�f�s]�$�!d�"��c�/���(ry�;Ah�ɛ��1;���4�����M�r������قm��~A��u]�Ut$)@�f�N�h	�>�+㼕�5�+'�0pԁ����pґ':\4�Q��y�/�<Q�/jqق��T���m:n,��Ў��u�v�����n��	ՊmO�/t�������)rƧ�
�ht�sq�}M��y����F����O3����`�>�z+`�_��99ԁ��)]�`AD�/GּT#��ŖpM�qY5nM��1���d�1?�H@{Ŭ����N�}W)�u��DMczo7r�����S/�F<(�a�4`�E����X����+s��3C�A�;y��E�SF|�p��&��[k��5�
]��`4���z^����u�gz�'''m7agb�)��B,��|�����w���MxZ�qž�ҩkq`fh�H�c����v��V��7<d�=�=e����[@��%r��	���MoD4����*����*��7\�\� z��q7�V�w�m 	`��(�5oS��5EI�w႗T�7ѿ>���y=�	���L-2����D�a����G���d�U}��T���3��Pj�S�ˑ���j�7���K�2R���� ���x��U"76ۀ$o�>MKL����R݅DT�M����ւ퓾��/d�阝:m��*�Z�������������DAr��5.Ţ~"��:-eT4�uIu�(�ꫧ��2<wͤ�k�G��ѝ�د�^�����vt��G�9\���7I��ˑ��b� �݀�d
��h5��A����VV�}��
v7�� �Bt�O]�H���s���%:U$����n@E2�Er��I��srND��R�7N��k����7�Zo�l����\b�y�`�&��S��qʜ��6�]��X�)��@=/��ӳ����&�Z=\��?�
伡����e���{@��������{��D%j�p3��E R6FE���n�RJ:��F�@�����E��@�ɬOz.VXI^����w�f}ʴ��BQ0����������!#�Wf��A��@[\{m�I���&�A��C��� 1}��2����w�Ze>��0��nC)R����a(�GK�ÝƊ`C����<�Pt�-Ù()ɡq$M����P��7U!��T���pJ�įk,�)���2��V�@��i(+_ǰsz�'�G%�����w�Dө�%I�iv�Z}r|.�kJ�U��o�֙wa���d��ica���8��꒩�*�P�b�9�:��?+?z���c�D<�q>�/a��l�yPK��{y�c^�%�����l�� xy�M�� R5i�TI��}�����*߼�3|0� �]��3�7�Ę�r4���5<u��#��Ĩ坦�ڸs�7�W|,�lh�8]>>����X�L7�I��ar�y�+�7�CUK^V�� �3��^q2 �-L��<�\���fF��Vn;�\r|jh���6��$n���WD7D�JK��.=�4	Q�'���f�������}p��ǈ1���$-Հ��;���Ζ�,�o�=F5>4�������m(��!}�p���X�*4���K�"w�F�qdP�V����D�X�����zF���N>�m�sk&ͺv3a7-��W�Y�keQО+L93���Su7=|�e�kp�T��*�_�6��h��%���.�ˊ�~��Ū��d������n��W��Lv?��D����:�F������I8��0�<r$Hi�a&�ޞ?�N՘Ajޥ��&lu��n�8nd�g@
����������y�
;�����N�хhD�`�!�ظի��)���[��kKv�$�A������혌CpuM�>������p��5� ��И$'R!�p�TvKE��D�E3�q�z_�x�'/�%wdW�0e-p����{7���������I�-�C��FB�'����G�l�elрW䍶zS!e�7�����a%��w�:��������Jv/)w�]T����J�H*"�wiU������',��ԡ�j����0���
\g�:�=zhG���(����j`a�k�Lq�����^pT��"��)�D��ո
*����s(�1�p���_z ��z�Z���=���\���3�΄R��=��x�:~Oi�1���1�_^e���IJ4g{2냱d�#_�t�����5������Wd:��%�(:q������mS�%�J�wi�]/�A9���Y��d^��{��1h�37�'HV����>+RnjW�(�	��p!`
������KV.c!�LA�}�S��]¢����'����T\8Ѹ�~��] _�z�	ډꍜ��`�O��K�be����g,1��sI9�r��Lf"^|�c~]tt�9b�B���;6h�,\c�M�V�`�u�!+bjxw�Djd�V4�*�#>ܡ�\E)L�	l��9�hȝ�W���!|������#��OaC,3c)�U�݊�3|S��57phG.�{B�?�uSu�۽14��RQ�.F���uP�+�:���\d�]R���O��|�\*�M)|�b�V� _A��bU�ˡ��{-�i�t�"��5�:Ib�u��Nk7&��U��L�N��$!�ږ����]m&�ѳ�9��|o�(��9��u�D��[��y�rY���.KQ���;zHCغ=�*|H
�+�^��KbG�}�����Q�aw1tҗ��c�P�>y���-$�Ow:V�ʷ��{�k}]�J"����cfeݴh�@ .4\����)No��0���-��/��Y)����0X�ҕ�.w��T2��D)"�P��_����.&�j��#R�䏰I
��hC�
������s�o���qhR]o�B��b�p�p5t��B�#B�u�"'�c��]�����"��:3�o����'O@'#��>��}!4��V��X�Yޑ7@ŇV� Ys����Q�mdP���C1�l����o�a��~����>��.���O�Ym�������m�+���O�l&��=Wc	��e곊��jq��P�k��Av��Ϛ2����(|� �{_��	3	��{׬E�_� ����	�Rf��������k��9���ޭ� .�A� l1����y�`�R��F��[0�=��ɉ���ON�x�XK���l�����g��)q�7J���6S:h�qZ���[v����XhF�'܎��/�\?��e�V���-�3�:�v�`�E�L.j��+����PW��.B��)^m>-4{�ܱnf�-����Q�UV	��d�<���Y務|yⴤ�#�Uàߢ%�D%�����Kj��G��!xa�B����&�k��R�^DL�pX��q���3�h�*�7nB$������j�֕m��x��������"�
d+'���(�K�j����f]��|!:�8�6E���ѩH�Ed�N6�����j������I��W�7Tj��d�|���v)���s&&r�������$����H��A�9�)c�����`�,�0U�JN�O���>����5��:5�Յ��Ͽ�~��m�ĕCg=C���!+X�.ر��=�|�Ta`�B�Ֆ�\�M���[n��Bb���5�ZBl����&��[��kVI����]���D�l���[6=�/��6N�M���5� �@����=O�QV/ /b#�2?�֎��j�����3�n��l�?w���j3�+Q���(3Z�JEF�7���t����[��u-9>��	��J��x�hOM+�I{#\��	)X��'?h����<�̦�;�%�ɼ�;�/�K��&�Yť�*��K�{���̾"	?i� &��n�Q��xu�&���<�6A�_��g�d��"���˧k`+�	�F9��+J��W"��Zd?�t��{���ʇ�-O)�B[�o�������#����i���c���ґw���t*�wUZ�Z����Z�HW<�6�.?�<� ���&,9���\�A
�Ӎe�'j��1Oq���Z����'��s�2|`V�
��j	�Ǒ�ݿK�K���2�Z��������d���R
ߚq�R�~h�@�L��U�hg9BԪ����yؤN�=ee^�Vyw��!��1��y������h���qD�Q�c�z&��Ѯde�?�[�(j�\�+��æ] �6�Y��%l�qG �X��to��!�US�e�n�*..58�	Υn�߂�n�X�����+sO��	��%���7�D��Y�"�v�0��@oO�&��0���(aG��5}a�ʗ2MC�_�89�'+QerS�{Z���GT�bw+[M�
�����(c[���	u�6Ȅ�iŉiͫQ�\��!�ˇ�bN�S�¢���m�)�9vj_�q�nK�������.^F��.y����k%�a�U?��@['�{��n!�2��>�K	�ن"*��Ɉ[�J�
銝qh�T¢���v/��x�!|���i
8k֎�i�$��CΈ�7��j�<�XG�M��LMí�xG!�^X��>�A��}x�{7>�� ��΂�Vj��R��S=���-B3ZZ6�Wg�T�y�*n �/��k�CCڵ	>��q���WdD��v����kD��E\r���M�u/�׶b�U�������~i,����)�:6ḭd��~B��(5�4��7�����f�@��7����f�Q#1R��&�A����ŮiԄd&���T��!�7�	��yo��զv���Sߨ�)FU�ahz~p�7[S���e6��i0�%�H���7Չ�M&��p�a�Q��RH8g
���N2����Fj�#9�2����
'pLĚ���C�zI�%�
ߔu���:�Z곧��f<i�C�'��BŸ�;�� �����7#O�ݼ�����$fU5dl�NO*Ύ�B�2��2������v���! 6Z�GT1�xtϢό�'-��n\mAk��ja'�D�ڷp�=Y�2ѿ����Q`��I7AV���hs�2t.�C���J��C ��.�޲Q�h��\z�'E�,'C��#���_S7�y�����j���i3�X�W�i��yP���	,�D���M�v��I��r&2#t1���/Bw�2eD��/k����=���S:�QEݔ���;hҊ�,_��ե%�'9��j�M�!BP�;b�(�'ְB��Ը�R5����UL֩<4fA�6�x��E��W�����&��SN�]g�m���ϞZ�����]�bw��OJRhQ)�`�Im�Oۋ|;�[��;����@���Z4����)Ʌ �	���6�AXlxVHYEB    4f27     d40%�`~��N�U��ΫӈRny� w���c�C��=5�n\9v�Ix9���]3�iB��q�~��5PzOO5����{8)6��#.ظe+�.�F���j�y���W���Ai�%+=D�'���05$3~=��Ƶ�Mm��7�}��ǭ85�܎�l���
1�=o���`ǐ�m"����o���9ՊbWJ������mjFN�J2�`A+�v�?h�c����q���t D	ጊ����k]�ȬsyXT�yn�T��utjoB�x�� Y���� ��w�
��U��-��~�&�	R�!�$�������؎X�LX5Hb'�
"���{Ӭ�z�vR���D�s�����X�C��]��?/�?�c+�\m�|�c-�y�V�F�\HG����Ew��1'Ԟڪ��Ǻؤ�3.Z�ĵ�ձL�Gn�;&]$���_,O���8*�~y����0�.n�0/A�۷�7�n󿹙136�PP\�H���pս�é׷%XH_��1:ȋKV=�Nն�	
)���T�PE��x�<��l��Ar�(Z����b�3���)�@,z��l^=�4��c)tt���9S0B	mH�������.O
���f�q5mR։;�v�wlx�%�,��{�f����D9E�Ǘ_V�t h�Y��ݓFI-j=��K��m�����w��f?u(w5Z�U�N�~1xN|��S?�b��,T#�<;`���<'�՛=yF�X��t:K�n��1,ڎ��Ah#J���m�~�)�_:[.F��\�٬�O�g�ك�?u�V}��ؒ�`9C燕.>�J����q��]$�.���^(���Ѽ��I�5�ɠ��#dߎx����V�'��Pg��X�H#V��@Q
dȃy������>흓l\$�v���[��Ր�.&�0o�����ɭ�qJRt�ni��M�ӎ�m1:P�]�џO�7hg�����x!C̚7��t5�[|P����a7�h�Q��h�ɗ?\��ت[�`¸]��ҏ�D�9 mJ�<�O$��n��Y�j�7�&�m�����쪫u�/����� 85W+�#'1H7�T�ߜ��Ǯ�$�?;&rm=�{�Һtg<�3�ݯ� >���>�@f`��y/��G��s�����C�'�^R�v��  �8ǟ����\�F�;����3�P&�+�ҒxMMq���Y�0����B�@��t�W�"FD;� @,S�4��� ɻ}}`��+���Fg�LeB�a:�PEP�!y[�T9���S��R�>�$�`��'�ڰ���g��`^��X�ia��x���q���2�3e��{�!�����$��#_���5����tn� Z��V��F�8u��3�A6�xl���* �_�=1Z�g'�8��~��$y��ds<}��k���D�F�
>����f�8�T��p�����X�+@zU�j&�IQ0�c.&�VIf�w���V��Ҡ�8��,3��r�S܄����i���vB��l��O�x��~ 1}p���E���/Y�_���ep
V�a:.0��`�(�ty��%?��0wݬ,�+9L�]@�$�ext�7;F^��u~n����`��H�q7��c�;|�k.4f6��εe��4���1WM`���Q���~\kW�Dt�����9n�6�Z@�@ح�(���|�Ze�$�J�59Hb�b�:L�'��	��6��Ś�\j2!�7URu�̭%�Ԝ�Ē��$�T���k�ނӆ Z<��h�h�;�*j@�G:�ϛc��b�΀m`$Ș���?18l]�9a�����?�<�a:�B�i��Mz�W�Ք��ybz�}�U��Vl�v�ڢ�i��͓���5��ă&��e���| 4A��&ʖҤ��P�� �Ъ�"�'լ����(�Ҏ�����X��53[���l���0d	I����5
'A2��1T*F�O�V�J��F��Qy�����6uUp���z���ZN7:���k"t���ķ\ޞ������.��LW�@��>�>�Q�÷�r[Y˭^�	�����=j���3�EO���)�
s���g�P�	G=�k*N\w�L!!���D�g���_�*��m�%<As:3ŀ�+���HPU�<� w���T�%��S5����u5}��")�|CeHJ��z�ﾡ�����3��똩����a��T�C��
����Idli��DUa�a���e��g��^8��4�����rD��͸�6rh�_��a�_� ���޸M���	)?[?��5�m:kD�͏]���K��Q�ziN[._ʭ��{��j3���v���r��0�}X-E<��Y�6AU�h�Cc�^�ź��Y�"Y*w.^|��^To��fΥ���Oʍ$�n�;,lF�I�B�8��7/!Buw�Ø@��	�]��u���.p�
�������WD$ѱy�&_D��dxF�u8��
05?g(	T��C��՞�F+�P���������H��%|1=�+�#���,����t`똰)��m�e����T��ԑ]�%C0�ɾ�4|K��}��4������}��*�|.���w��u���dc��O���#1�Ѓ�\���g�
U�B�r��^��D�K
+(^�(��b�$=Q�Sdˠ��`����a� �A��1J��pe��:�<��x�+�tы�uG��N*0������e����á�� 0�h�3Sr� 33:r���-��Ǟ�v��@�T-j��!����D8�b�vڰX�f9�A��?����mN����wu�x��b��T�n�\�A����%���:�qI1�m`Q��,S������A�a�HaV���Yt�N���GUR�ɵ���۷��li��I$�	gN�WY���Q���>���od񲹖��VƼ���?AB��0
F��>|�S�d{Ջ|j�a)���J�9���� �ؒ�]�7P�WhX�|�I�c/����C?��;�M5�Zs��N��5�_��>`�A��3���"=OŅ��a���ӉwrA��O�\�[^y���)MJ��a�)�uY�7t�2-;�}���c��uPS�MCyʞA7�Q�D��Ӡs6ѝ��B�C�����`�'�+�����S-���˙�Ե�n/���BtaI�ΩT��1a&&v�r�V����YBN�yo\|�؂m�����9C��1z�������nΒ��g���_�}|����Y���T�1T�Y�}\��뼪��M�O�;��2�z����N��������°X2�l�4�7��Dd�VQ��8\l��x�)XK��,6�?F#\6J
�LL�=�'xX�,g�v��{�}��	&!(�^}�v��e�Cd�