XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@5шwg��r��/9��{_/���Q�A�m�!�7���̍��D�kӧa�JU�f&��a��4�
�dG{v�q�dH��m��Anzw8�?��?x� ���*1蟞��Y�U�8}��BC~��&��~�0���\:�R�\}pV2�B�^�_�y��z�q^����@|��td)�^=���q&�G��0[��q]ZF���7f�.��N��K�`xs9��&p�������0�!�����T��x����@��C�7jC���c)�K&���?P�B�����l�4Y�TL/+��e���DFG]~ϖ�����?4�D�'X��h�	�b��P���;��HJ��y��F�E��Y�=x�
���F#�e�-���G��F�֨��JM�xw������sτ/m�Щ�͈�t��	yM�K`�?��'�a�l^6���T��v�x�+`!Ǻ|��P:v �7�wUmv���vý��(ш�^0j���9����g����Me%��'����R]�T�M���X4ɦy�c[�����jO����iRĐ���h8��*z�#ؾ��|�P�����2�x<%��o��[l�!@3�w�w=jP�p�$�Lr�e�����*&��y�#�B|V~��{�E�m#ncs~�8C�՝��9J^	+W	}���7FL0_T �d�}��T��Bݝ��J����V�?���:ZJ+�|�	�-+�1�3��\'�=T�|F&7fp4��E�N�5�Q'�������8�XlxVHYEB    3b6c     e50is,-�/�% g��3!%��0/�>���2���>B+�h�V�˳��o�/��z-��������D��JY�yf6�հJd2�|4��T)d#�smVb�)���xŌ���sK_��P03��+�)��ME��ڑj�fL� ��ֶ�ȑ�E���9�
���پ}-u�2��G�y�s�'�࿎�?��y��jZ�����^�ĥ<�N���N����L/A( {[IV�US͒�Ö�z�$O9�o��o��S�6��H��vu�VA6��5���GU�H��6�>u�:�iԚ2��|3k�����ErB��$\��}c\��w\��|�Ѓ�	H�c�<���I��l�&ZB6m��;-������6�ۈ�!O�9�(��Gx�����/Ə�l�ޣ�BJ�Q�C��*P�?�4G�22�|�|mN�vGO[���1Y�Ё3�.����&j��ujS�]m�D����i��J�\Ɉ�{/:��1^)&Xp0��lT��M�Y�9
@kg��'6W�8&)�:��w�����B�xg�fI��;�H���K�4_J1���X�o^c���?��+�����1^�fA��4�آ����Xf=�_�ӖrB3���~I*�G�L����2����qD�Yl�O��	頋�0W����N$
[���V/C�5���Bv����v0H�(8�:�`gO6
��f��4���oq�j�7���n\{�ğw�2��k��#v Op�����B��?��0��i s
X��#]`ವ4*�-�Ʉ*����G���[�VQ���&0b��i�� ��]:�\tv|�.v��z�M�M���6�s��	�/q��>���l���)��V:�t����krr o���� sx�j��b�3�S�He�������������G�d}c����p�J���h�4 �`[�"�,�z������������MQ�#Ss�V��VH���v�#C�������~�4H�㗶��������u_z%dC����a��J�����5��b�.�hv�Zdk��3�!���ȏ*�<1�Z�U��_!���M�B�����A�����S`gw�G_��k�h�Y�ߏf�l�P�h�I�Ia�Ҩ���n��J�f��-��`�N��nیa|g+{��~� ��*s*PE0(�Pֱ���/x��s���OÝ��]�-H��I�1�jG��Q=�Y��N��ׁf�n`Wa�C�]�iuwz�b�,T�LWxֿ�ޜ�1�T��Ew�KTqjWW�j�L�p�Ũ�?q��X��lL�n��^q韸��u�329�nK`<`o�A�a��s�S�N��+UT�9�SA�i#��� �=�Z7�W���z�B��?ׇMz h���5�zrⓊ�?]yN;�d|^V"��L���+|�&9�5��z��ȇ��N�!FU�Xl�:⃑;�9?�~�5�6��"vofY<��=����q/"�$j�< >,��h �ig-]��i�Z"�ť5�̕��A�=�\���y��Z=���������=����K�Te+��F8��,����6��=b����G&=1�İ��.���K�t=��槄��i���9[���tUhqa�F�����I�u7��*Mg��S�%L�1����F����B/9Z�#�F�{���B!���Z�����q�";����:>)��׶F�I7���L�{���Y{�2�D��Y'�#����t\Tx�p��w��
,w3q_w��@� �ċR%�/M|Y2�����1�X�xPЋ;�6�l\�0�j��KO(�;�U�p��{��M;D�^<��C�lM�?g}.D��12٥���$@W���P�l���]{�
�1��u�I&���h�ҝ�1K����xu��}<�xY���sr��C׭�����<����+P�l�F%£U1�|�`b,�)=%Q{�� v>�$]-]��Q#A7��O�m�)� ^7�#�����T;GD����ڙ��^?j�A)gw�2§�Aع�����T�>��r�q!h��Ӆ&>�tn��C��Z(�Eq����bY@H?������\��-���W����,0�;jT��Y�+�:k��L�`-\��
oqñ�n���Y�o� ���.0�Xe��1
�A��f�4.�Ǩ�3�*��UD�~X�>v�X
�=S�a�4�5tI�9%k����Z�B�"��Tt5m��..Ҝ��Z�(+�BmU���OLB��'9���y��_� \�W�j���������V�;26uݦٷ]��7�>*�h����۹�1	ơ����Co��Ĳ�_dJSG�K�N�ΈS�;T�[� ��p��Ȧ�x��s�3�pP#Z�T]HB��NѰ7H4*���A�G�� �?�]�NHyGƺ�i��Y�\dN�����!��S6�`�4�����L)
����m�R!)����ND�$�Di'�����?�Oa@���B+(��KzP��N��mc?�挆�C���'��^E���~4~���W�5UT$K~p@���GW^s9�Qx�D�N��h=G��T�CY�r�:zao
͗m�EG
jrI�Y�{_�~c�s1݋_@��Rq۟�m��k���&k���~�����7҂�n����rB�Pݘ�J���h���`;,w�S-���c�����9-8�1HY�ްW,X2�L$gb��Q��7��RZ�@˗��j� ��?�RWpmvၜ�I��4��55�_\��c�D%��8�º��E�����]��w����K��Gv����\�L�(%דyn������� ܟ �9Kn��ɏj�xD����*
��oU��|�qw����t��嶜�{���I2���J��@ba���QjVW���9E���+�2������c���+��S�k%��~Q�0� �_#}�\o1�Vq�dP�h�������� �w8n��0s%@E���^-�!%x'�䞙3�-x� �q~�h6K]�G���?|�[V �M� ,s��.��# Dԕ�O�đ�n�-��w}u<6=a�7RͶTl�1eZ����N�S���e���4֠7 2�z��b��Bu:�=�r�2�
���q���.��w�o����@Ѩ��Z��r;AZ9v���h�տq�j
�ݔe'g�"��x
ΑG����	#x/�d��oEK��>^?�_x�\"���3���@��É���8���5W��;�̛s%M��ںyyu�J��T���K�ި�}°ɭBvC{�f9F�Y��*���۽�a����Ҭ�"6���y��Bk<�6��,��0eR���@���`�@�P�o�[ ȕޯ�WB���el}�?�]��+�hB$�ŗ$��R���<~�*[I������"��ȡ���G�+B�d����$�� oʯ�3�/B�BW嵍�,-��g��]ց���%�Q�
���l���@F/+V���4F���������E�����������uu>�P�)��o_�b�_K���-�X��[�?�E#t�*%�v>��H���v���-�`QO��]��1�.�UϾ���K"	H_��J�H	�6��&m��&���$��B