XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m��ͨ��A�`g����i8	:��=�+^n��^i5d�*j"w���v�RP�P@d�R�`,
��w݀�Fb}n�Xk)��K˦��"�3�KW\4˕cqHI�#%�u�|��mn���P΃�l��Z���1�\g��8�����=�?�qzܣ�D�س8M��Λ�TH����͉��uٳ��}��f*���~�UZI��8�&�gl��߲���X�-/7��+��!���B����8�v���E���jt�b>r���8���	揨S��\�\�H}�D�X*A��6�nnZŜ"}�}��̇�èa��b�vwP��>Z `)��I����[�zo�)eiV�������R[p�+0h�E5���!�s`��7�4�G줨�*�oJ��%�R1'Ǩ�`�J�n��L���c^R\��=BEg��䥵���A��Lo����X Bf���K����[( <�j��!9b�<����u:�=�h� �]�!α�b�+|�T�N`Oz�M��h�!��R%��i)�Տ�o��N��B�����+�)RD>q���5�W��!��[ct�{w�jvSV]��F�_b��w?�|)4�ٮ;��?���wY:}��n!�i!wG�%��� �WT��Ȅ��渄c��Ư''j� Ng�"�OJ�Ǐ�e���, 2���]��D��qD�$��K�#��������Y�$��!�d�DQXQ�f�2H�R��	�AX�b�D�*�;=���5�]�ĥ�'�%\q�D��XlxVHYEB    117a     710�����.Vߜ�8�����c�&\�צ�ָ�7�+9Jn������HB��_�a���/⺻p���?��g4���4E�P��Ύ'T%��{"��Ϭ��k�:+?Bʾ�ĠV0��y�����ff_-��9qI����?���e��F�<΋Ý6:�
 ;�9�T�e��Ѵ`��n��n���7�#HE?������Ī�|NZ��ڛ
eF� ��φG��`jl�Jŵ�9埻��=��)K>�Gb�x��G:a��te5�v*g0���].���S������x��i�[�&:��R�Hϛ����]�k�K������.8��3��f����rHݝ�8x�d	n�Ú$?�y�l0�j���ZR"c�H���MGq��K �1�4J������ٔIݲ���z�1>�.Dʖ�Ls�����=��	�Si
��W�PS�8=�����n�Q���o�y�S���6L�`YoYe�s#T��o��`�^��	�.|�X����3�D��z�jǄ�>�0z����a�X!p6x�-�Z��Ң��J�R�B�i�-bx�����QF�e�9!$:�+ޫ��� --�!��=���+���n�5z�ED�22Q.}2���;� ��z�R�2����.r]�z����S��<F���Oa���)[�7Tm����F�~�Լ��t�&��Ie�?��o{��16�	Fs� ;��^��Mţ�4��jB��0D����!�,^��"�:�h�󂥖�F�x��'��KV[)��jS��-�;�0W�#���<�	@�{{B�
��6Cߐ�<cǷ̈́��5&W'��9��fH� �(��1�\hr�
��۸5D�������1����0H�	?IQ����uL�lg=G�n�n�d�l���2[�@-ĥw)���x���k=���s��ЂM:S#��c�KWhI��G7��3.��e�z���\��,�nB.���V�RN04��N�~��A
:��i]��eO�2�X��XV*X&=t��G~�Nu� jd�㾿��ٷ:i�]g7�s��C/(�����>w�}	R>)x�1�cf�A�^<#�&KY��)�.��D!>�|A����>)�aro��;��e�P�u�X����y��YvT��Š�ΒTK��5��D���Qظ�+Y��E:�|Hn���x*Y\J/�����B��0�1{t�q`��ʻ����+RR2�h�u�7 �l��CPRKR�������v{�	=�9�Ն�
�*}���u��fz�@��-���|p��H!�G�E�������|�����ŝ�S�o�b��l�G|����
������KvgOm���U��&'���qa�JY�H�8u���%+�P��H���3���!q��'w]y�ܒ
q���3�i6���Z��y.�1�f�;��s�"_���V�u)oz��H��j�Pb OiU�aD����`4�K��F��ёh#b&�q+ja�������Ú"mN�"���0@���.�YJ�1	�`�Ԣ�O���#����!|'�c���C�� �Y�������-<=�ׂX~��6�Ŏ���4h
��I�������8�?��HUN���ט�r:�X���,U��	8y��k](>��O��@R_��� ҈�c�r7���&�:��~oA��Q�tgEa�%"8A߸��ɒ��Y�YC��gR6�vΛ4c�@'�I����o�5ur# ی���f��ڹ0`~��P`���mW?�lx�K���꼁��J��9}D��&�-�R:��,D��U���W%���-GZU�9[�����N[�"��^:k���