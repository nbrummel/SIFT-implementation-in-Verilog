XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*`2�<1�n�������3�oM9��I�q�/�Vݍ/3�|���+P5��!�)�Cm�mS�m���n{��F\JoCu�w~���_�r6-!�4�a� ��v���l�Rxp�s�7D���)5x˾�U��
^D�#8K�`d'r��z�Bɔ3"W���[z-��N��^�-O�zJS�h{�m���7%�����������2�����F��1S���[|X��Q�����B�hu����H�\���]?u����@ �*t�iA|���H��Q�gc=O�B� ���k
:�6�Jc�9��#��?ꬑ���HZ;�S����=�Ֆ�.X�&�<(���^�Vu�G�%.���	|���qi�f���R=S�К1��v�,� G�2*n��b�u)�F��T/��a�uժ���r��� �tW�i����|���@��Ɩ/���o$�4�p��Vc,�s�!�R�><�������d��|n��_�!l.��+Xx�2��`̽��Bkc�*�agh�v+��6Mrc��61�\����o5D@�3�[7|�P,r_�I���͞�r�:G�X���q`���A�a�f�@��k���"K��	(�+=��mC�����*����hϲܕ� ��5�D��Pķ_-�
��.΂�ħ�3�<9�R�����a���t%!�օf�,�Uw�ʓ��g(��N��Ν�J�/6ސs�C����՗$Y�+��G��:�(^`Ł�8����v��BI�8%��jAF�޹��c:��v��&XlxVHYEB    20a9     a60Q�7�׶�a�db�_�E�Y
�u��FG�<dFz�G�'������'f��Bc����(�N�i��k=cC�Ⱦ�^��2��Ϯ0��?�:�w&Mx�I.~X����L���˩���4� 5H����B��`:���>�яW7�gxN�]q��+���$)�����cA
t�B}�U�h)���2$b�ZH;�y��#��b�j��PƸR�Ȯh�6�dUx��Sbd!u��@sL�~��WZ/����؝��@t�Ջ��Q�g���$��s��j��d�@T�f�'�%�ڞ. �eR��Pa�ʡ�̡2�Xd����ϔ)�,`�9$���w�~�C��䱤�&����`O��q4a���#�DX;�,���G� ��tӋs��X�8�"��?����N������<Z"���87�B��Q�(4�S�ҿ��ݣ��6}�G��ֻ�}��U��tm��+�^{� �w"(�����������)�ޏ|^F`�a)Z簦�QO#�����M�B��-f��3�þ��P)��c_���7_�X��t���ȃ�%�Fx�X�ؖ���a"���|�2���p!w�|�*CRb�� �{��iB͒�S`jdn	xFgu9����"7��o�u��m�U^0i��S��̟"�0��z1���A�gވH�`�Q�v�9��Sb��.P����"��Dc5u��>� ����i@ЕT�G���{#׵�O��,?nf�k�'.�mD��y���}	M�U��&/(�� o��w�[ǘI�:�4���R������ ?��<ryB�d�w�o�E&�����5�Q�t��l�*8v2ַ*�ÑEB�]ڌw��sJ��ns�00Q�j7���qF�v���]�Z}t��A�e.�ՋȺMh�6���ca���b��2t`��ryI�*��F��c�`���dB�~����5�$=�Զ�+ƣ����3�P���1Zx���:���f�?���D-D�	&�rЦ �KQ�6��є-��{x� ��&�u�����+�ox}p6;�5$ D�Rܧ4n��<@R��VQ˙�(�s�>/s�&z߬�{��ǪC�V����bm���(�*�أv#M.��_�<m��oI��Xґ�8�_JԞ!��KJ�\Exw��Y�,���� E����v�dizWo�<�X��2�B�2�p�R)��M�O
�'��Xx&��1���Rɑ��JNL˒0&*�V�fK2#��D��w�F�O��5��7o��s]w&��2�f���.��&��*;�B�m�z*G%�kØ�դ���R�! �K-��-C_�_V��Cu(%�­c,M�:�7�{ᛏ�u���� eջ�rJcg�-\���m(C�6����A����>�
���
��e*�*�d����-��XW���S�����׼���qQ:B�tw!�Q�����*dL���>�y{�0�1���8v�2�Z�C�͜ǣ�Ļ�M�HD9�[�b����X����F��0>b�~�Z�J���2,�U�F�3ں�D�3��֩�v���nȺ�+�΄��G�W�ٟ�^d�۬.���*+/��qR.�[�k��q^�#}Gv�:��� �re,/�R��T!�u���;سH�McQ�mڴc����@��*�_/��ZMЂ�kzU���� ͖ĺ]CߔFϾG��{��%d��7%]ƪ5� _�B��E;Wq���1o˾�}R�'�H}���Pv�^l>n�ѡ�& k{�$N�Ю0}���GǩqI��}��*l�*ٚ�ԝ�GW`���	���}D�K�P��^R���L������:]��?�,�ҡ7�����!ZC�{�{Aj���b�=3�xTK�]��J̷C�[�?����I�����b��v3O���pWU�z�$P��7�i!���JE;"�\��]�6l3:1���R��),3�o]����n呴�j����Ɲ8���2���G���Iv�
��Λs@��Q�9ə���~.:���D�Vb���y"0�A9Yn�5��3I�9�pt��b�n�٦�F�s�7���B������46<��z��-��NP����fϰ_`�`���I�ւO#eXy�^���HA��=��BF�p}�d�D�d�����(���+��[�=�����ݑ��x�h�b)��~�O!G����� _��w��!L���攱6��w����^��N���9��
���E�C7m����.������i�P��I�w�V�����j�A/W� ���(D�����^�6=�¿�j���i@����PP{�]��O@�����{Ujq ��,�T��gw�a�de"���)�":d�r� ���
�b_������tWvd�c~=�����W �͗���e�ם��e��Ȗ��Ur�B��j�w�_y���8�~H�}V��P7��f"�^�gӞ /'��a���t�ep�ܱ�@��Ԭ	���{v����(I�K��s�r�4���A����S����Xf2+r�g|��r�����}�/㯇]�Y����X�R��/DdR�>
+K���:�z�d�p��L�uam�6F��Q�������y}`?�:�?�D3+�<�M