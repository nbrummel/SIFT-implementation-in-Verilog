XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;����mrJ�w2�	�}I�p����˷���<�js�����cN�w̌ǟ|�t��Gֻ�Ę��k�t�^��I��e������p�6�aـ}������^] @�����_��n��E��vq���;��r�����:BmЇ�P��[ԶX���{=4���u�Ƥ�C�h,m!���~�6�l@~�C�y��7R��<a�����������!k��[@��u�I`�@�E�0�Sv�Z�G�x�Wї5���Fĉ�;j�8(m4�9�ĺ��U�Z�3��GK��]GP���������5/�b�6��gLV>��Wr�xs��O�Bv <�'��T�c+�n�-n�v�U�C�^����CGա�G���^l��*PA��|z��m�3O�����tbu��uL�B�a��'�2�=��?��,�p�al�N	ʲh�t�f�RA$�4��h˻��J�����9�-���`��\��E��ǺfB�@�&�X�P$��7U�]�V��똨4[�(�*�H���}����{��Ig@���n��J
~����N���@4�_���G�n.g��l�b�l�W�|*�cλ�ꍳ)���g�m�폆:#��_��0i�Ō+^�S����c�:@m0'ߦ��󷉊5j��)}�j�#����	�>��j�r����*�'ؚo�C�ic�x+����ݪ�)����'�1�^q�d߶ށR�cY	������X��*`R�o��^R�Cb���������^XlxVHYEB    4f43     f90��6��c��T<�}��{�_�}�D~���ڤ��<_^�1�,�8\����R��o�ra����5z������5s<>�����4^�����;*đ��8Wc/��m�a�ҍ4${�NK���#�'�N��@7M���ɣ]M0���U�b�}�=uu�RO`AO.ô/'��	�^�YN��	#�߭px4!�����A�4�%Կ�b$^� (���hk�+F)��e��z�}D���0�]X��'�W��4ŔڛqX��4�lA5�Drڊ��vW�70�\�<��ܮ��OOL�3cTㄶ����.��[]� 02�������Ҍ@����}&���0�	o��Ƙ�mV9�,�E¾/�D�U&1 ��W��4{q'(C2��=Oن���>�����1�I>g�׉��|�76�Ȥ���R��r�����A��y����L}u��z��zP�үhU?�ؓ�}�A�ł͕VQ�x��|�0����p�G�&�v����D��9�س���`�+�(c�y�)��Y�(ب���I�������J$5�����8:'k�t��ut9�noq�9�3���r���^&���k���YKC�;R�E��.��6kz|Ͳ��I5�H���%�e�K�<����/9c�)�0��?$�D��qg����%>˴�<*N�h�ZV��^��]s��]}��[��<x[>�?�N����c����!Z�)�x.����c5j�jO�,߆��+o���mf7Zrް8�����̑{*�W���M����I���(={���x]ّDW5�r$��{��F�v���2jnnM��d��ɘ��	�q�7��p�XX��n)�a�	Q�����x}���<R��5"N�hh�\`��kU8������L���w�B�v.�8������ ���nN����;cG`�����E��s���6d�w�C�j�����L-���&�aQ�|+��J��~{�*aO������K|���#�]���r'c[�����
z_4P �T��E�T�GQ�Lܢ!F���>m���'&�t�ȥv1�V��"4ݸ�$2�<)*T�����96�j�щ�5ԇ�H�[�bd�X>1�`]��M�O�P���Tl�L�Ye��{z2������]�b�w���~�ZD8�f"�
�|&������=U��r׍	P���������/����`|���� ��C�ſn��xh�s?��N��,���vD�h�ɖ��8����w:�dw6jگ3z0
�c�uGlS�<%�������Oج7���`�+r8�aKa8;���l�n�Vx���o�<fp��3�_�N��b�.�\VȖ�pS�V?;��,
��li��!'�1E2p��@hm^j�����X�S� �W)I�^*�X�ӚH�b�f'J�ګC.����"�뜷x��m��/h�pOW�`�~�G9g��c��׌�g}��^AF����V��QJ`��?�G�5�H{��ڈ�Ȋ�:��
Sq��ϖ����o���X����^.U��O��%44�va���~\�o
؊�� ��(b5��������ңc��� ����J7�U|����2�T��|jI˄�rn�՚o��=�Ь�Ǣ�?��T|VHIo4��� 1�]� ������%n�ѣuvۣ�?|J����Vs̷�\�*0TOJA*���=L+I�Bu��w�*��lQTݍ��Cbk\,�0G���{$��������7��#ʓ�we }G�_�cJ�k���_ȅP� 37k?�.��-R���	z��Ӽ�y���!A�.~�<dru�?�Pn�nݹ*�v|�fo�e�Nx� R���~ɅR7gu���c�ng���|=q��T%���"�ݸE���hƳv5��|����Y<�}`�G�`�]%�MZb�וk:�vAle�T�- �U������/,�B���	}�r�N��[�$��
� t�j?mHz;�$i�ʥS�olT���	Z��T�<�[���������U����08�hE��f4���B5Ǽ�1�Л��2+���e7s� �4�-r��P�'ru�cX�����"E��j���o�EA��O9�?���C��Ȃl�Q��뾩��L��!C�����qB��=-��!a{S} �R��B*][\���Y�)��+�B��gD
��-������pQ����N�����:��M5#5	�.��P��٠�$r�`��� �/�s�3X0>�B����F�q,c������xK*���&��%���$��i�o�][�\�-�x6��	����ůݥ���-v,���0�h�*���KJ.��;��=׻����@��qDC�Ǆ�I�
W�Tw3FJ��5Eꉼ�D�Ж�`����#�i����ޔ��	15���b�ox�m^X������;Ĕ����J��)��|�0;R��� Xo���C�:o����	�z�u�?qV� O��r�WVQX%н_�vI��	�5ah���])j�Q1��g�G�1�
kG�Eq��\�o���j.�p���o�8�܊�:"ƣ�F�hLc�J��-п'3�n+������<vRJ�qA.�<�O�*�^���8ʺE*�J��91��k44�x d�ā���7ƵA��}*2(��,Q�q��𯄕CN�B`�̬��m%�yJ��g��5{�h�c���[���3�v���`(������Ӱ� b":�N���ᦴb�UR]z��Ӓ5�����N�1?�T�A��I��?5�DK�8n��그d|3ޕ�����G����'Pat�I��\����5z�Ǔס���> ���j��Ys��;G�:=�
�.or�:|�_6J�1�D���f<��!��I���~�����ϞS��$&[�*~@
[٩�HM%�6ҷ���do�F����?{�����s�����~.��~xG�tNL���9�	���a��ɔhZ� ��"�>��/@3�,2�T�ΪI$�� y����q��� ,$1%�i���`>�(�,P�7�#�;���"���Э���ؑ�ˮr�sT��}̸�e���>S����m��\I�T��C�Q����W�[�{\צ�N���҇���?1(�$��ȴv<������}�:�}]ΌYM���y�����lMω}ܵ�
_c�{
[.G����WК0_ Ԏ�o���c744��J6��虎�+Q/�Ő���f���%��/
o*!���
d�c�1����!s0����&��sI��m�14�ř�N�Q�>n\�<�+d�T�מ�H N.۞˩�����`�
震{�^��acG�����lM)���S��p&`۷��	���o��4�ٗܧ������b�� ��8�ͨnt
?����% �!Mo�,$P+,���3�E�
�`���{�tD>�Q�v����\��J4����w�"��'�IY�����~�3<��Ё3�a)�=�P2�3���PCz�zئ�l�V�P��j���OQH�[�)�w���Yp�@x?�лu��Ҍ�E�d*K�L�$�a��$\�X�����x��$��a%+M6C�����7�b�,��<ǅ�a����T	�}<.�y�=N�M��/�/[�Ba��p�p&�@M�������y�m��7DE���c֮^B�������|���H1��2��k�E���a���qtI%5j�����T\?A����Ѥ�=nr�9����z��B(�X�#����VIn0��8?0��O�ؒV�����':fV���)��d���O��TU%�W����D��D*cW<��p($�L�h�o��0�?������}�8�|�,��թ�[%�L�[ׂ�qM�1����qS�#��y�X