XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,��˼���E�.��n������j��&K{�7u�@��x0(��RYg�q��@���e� ��Bf�e%N�>��A0L�}�n�+��X�N�*_��qfHlX���"�x�DTEn�y��(�[����W�
3�u�[#@t^�Gn��[K��㳝��^����?�ݲ����/�K�H�_`#�4��A��|^ϩIH��w�����
g6�9F;�Ы�<l�^�T���kuׇ�
�I�W�TO�I 7����
�YɌ��	�1�f���~�؉}�5l��w��d ���.���.����O+�T#��5m,:�c#�o0W�.����F���S�����7�b2��KSA|Xj���N��E��ٮ�*��@p|�TVY��gM��&�Ğ���,��(=����/��_U�z��(���l$�K��}���|�3#��b��>�%n!V��ΩF-J҃�et.G?GH���6���*�F�O� �
�O���Jx�	��h��6��=�څ^��Pa��Yc�Z���:p⺃��tx��>�a�o�����v����a�̊�������&�X �����Bm2��x�;�~�]8���P���2CUv��<6pi,�/`���˱g=l���c�z"�@3�_���dH��P@���"��������/��6�l7}>80lr<�]���ۃ�����&���,����X[;RF�#�jN�0�bG���G�X���=��S�/p.T�����c�N�ؽ\�8��� .MNU{M�XlxVHYEB    2533     b00�`�x�]M�Z�_�7O![ЏTV_(�ń��j_�Q��9(D�O�?4g9��𪰮�i���B�}��G4�#ß���!�v�:ͥ%���F���� ��Wr�(�;\�v7�浶Ɗ�����aڝ� �8�:2L٫�1#Ʃa%d�ȗwU��́ �f��ʳ�=�(��J`��.��	"Q;��?7[�t�xQXfw֧���ׅ���\Z��59�*#r�<��ފ�Ƙݱ*�8X����M멌�pV���j��"�jycP'��}ͷ�����! 1Ô4��_һ�Ӯ�2�HIn.K&+�-����Ě����jKhA3�%��SC3w�p�����k!j$֓dd��a�8$$�3E^�����N2��z�����L�f�t�g@������ݶ����r�C��z!E^V��'�,]�&��
As���)b�!pJ�g�}�����0�	���$.�dTUrW�7�YQ4CٮCIo-�0�l/��݄~.�*d�綪*so]?�mI��@�r@��}��K���P�Z3'R�k�
��3}��������
��s���Yi����(]�ԼɊ�˃�)R㭢�_k����P��E��@�!i�mɍ<P�oF{�=�>�tՐ6ų�踱p��n�${R�UǏۆ^F����!���EC� ���"�h���)/��Yl:�����*6qPuQ����ix�h�>�]~Rg`�`��ZZ����ǢT����]e�E��w5���D��t����m���=�8d�t-8K��6[�V4wum��|���,C�=Ge�Z�w������@��jg�Hk�u����O*8	�k�b
E�gŹ�QNL�a����{.;U��V{����\�\��g���'{�x��Tg��(��kI�%�F�tN�rx���Ȥd0LP�=੕�<0*<H�J����n�$j-h�'��k�^ T@+A!�%a��7��ܜL\1i�%'FcN}G&��fG,��9�A�=5�������w��`#���1K�fC��LB��H�� a'n$����l������E��)�!嬈����͂
�|1h@-�L���z��L�Â�ym�I�t=�g�k� ���O��j;oDꖈS�V΂8 ���5�����K0�DJGHBh�[R�0N%M�� '�4ݷ�߯�i�~�i�}�K62-k*��k�g*o�#���D��9<C`�5<�&�P{SXh=�Hz2ˬ�Q��p��M���MBb!���'srr[�A�&�L%�+6YnB����He�,aj�� =�{��K��Fw	�G�K����{�ڂ�������(��r	w��Ҟdf�N�1��!q���v�8�Mk�������	$֑쿁u�DƘ�"=|�z�J��z��+h0�|d��*
�(�-I��^��a�a�]/2$/��%��b^�x��@�������V�o���M)܁�&�[�_P�%��<.)�@��8�%��4��oeڵ�sr�]o��.�R�Rɗ̝N�UK�+�ZA1�����tpأSk����0t%��Y;My�Ѻ)��y���q��LjUQ�^�����RB�"%�a��S�����n�+�{�"T��f=�m�jzƔ����	��w���ީ��f�eOY04��́�7U�|B�&�%yKp3E%jp���F�v���d�$%.̔6��zb�C����Y?(r@ƅ�!�7��/n*W>��� �{].��	8�ZB�W�.�q6�TGimg�(�$� �����1�EQ߁Z'�P9����T�us3W_SK��.�D��s�s�_:���_2��l��1",�!��\�v�t�x�~�M�ə�3݌Wn��@~C�t�>%�f�.�oPB����ȿf�?N� �=X��.��(q�cN*��
�%p9������ `p��G�3}l$ĔZ��(O{�ɸ���38����>;�W%I��dY�n��}����.� �rW��J	����j���3V�i�QqO�)̨��ťp��5ﲱ��K3D�@�׾~,c����E�(I"8|��W@����Y����C:L�$x����&!�[c�.L�����D����FTJ�cD-���2�z�,���l�q�t-��}+,�a���e8~�j�-��oʓ��gp'�&*H���86kڬ��ov$��zB��w�p�P�������Vd��D�V�僄���I-�.>�=�;ŪfV�x���²m ��IO
()�יp63�-E�t$xR���*����T�5ڄ ��pv�t�-�/��h��@�8�{/���
Օ�c��q�� ��%�b���EeH��CᡀX=�(0���:����ֹhY�y� u�#>��A����D���X*��QF<���@�sC���P{]L���}��T��@�l䞔N�%�U�l�\�����q\��B�p���xB�m���h��y��ǖH)����e��r\�2j��p��1-�K$\�Mv���|��*�N����ڨ�#��O*����A���;�i5�UVl]ڢ��v�F����F��k��2��N��J���	�ao�P�-� �ë��:�	A�J}��:�' ��C����g�j���x���>2<��3��C U�q��)b����L��QW$ap�- �����	��]V�G��m��ѬD:D�!*�A�|���Jk�V���'���xj��:e08��eFL%4���B�Kʽu�?��Yf�J�o�?�����*�_�~a�2Im���H���x��Z����ԣ ��#$����\Tj2�u\��y��{�bg�w�J[�