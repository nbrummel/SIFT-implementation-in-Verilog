XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��EVǀ2}�����uH;�n�m�OB��@��E^<��~���p�X���)��o���xl]G��`�x-d=L<
8��#a���O�}�/i=:k����`uX��NR�C�\I�L�1�Q�\g��?:YӴ@v��R\�fM�_�'���~m�ح�[��m���ZK� �ZMKwxB�l���f%L�]�]w%țěCN] /��T_���Ǵ4ViI�ʃ���ӎS9�Y��>�����'<=�UgҺU�l�<�a
89v(��
��#����N�4-%�x��u2�AQ�����RU�0���6r7���:������R5U{k���oi~	8=j�W`�5��ӱH(rÌY4u����l_�����V�;�O+�U��bɑ:N���+[�dg���F�����|�w�$����e���n>e����4T�#9Y
���]xk�����o�����"��)�8�1N�ag��R��x�i���n�pcU������O���3z��X����@����!��g�D	�.�X6�g��m��� �.�x�xcۿ�:��=S��|�<�fdh'�S���R���S�m�%+��2�*
%�<f�4�y*ի���q�/�j�-��D��O��FX��m��gN�;��C�`��K���#7�{�~o�?!96��!Kf����ò�;}W��o;Tmv�d
~��Jt�22��D�I~#�8�Ye;�k��j/&�U1��xي.2ӌ���,8t���_��P��;?*9���<��3VXlxVHYEB    20bd     a50�-�<���O83b0
�ѦS�L�!mw]�m �p��"B��( ��85zd��D/SV�ī�C�膓W�~HOPXJ�T����eHX+qR'�����W&�I���y��/����Χ�C쯓MMɺAD��iZ,�rx�b����ͯ;���q�W��y�?\;?�Ē�KV��m.�򶐐��Ŝ�qB��'XSWTİ"�p��S���+΋��숺������Z�&&���+����e[�=7�ְ�����޹��
�f�U�_d��cs=5=m�����=,s.���fz~��ʢ ��v����[w�rD�5knK���mڑU�Q�3��7����+5����(຿S)A~ɇD�o\��8��S��B�Эv<����!x�L�]�Ds�vIc��tz������B�ig��{o	c��ܫ��2�<" �u2�B$>1�OyX>;ܶ�G҇�}�Ӟ���MF*���z^}t�����G�����j'�,y���n��Q��<q���?lyI��:	��J_��L��F�5����L-{�=�>�0���a�+
�.��j�a$�xw�:��` U�=ň��#�����f�X�f�Ve�;��m'\y��b����}uʅ�"���]q�I{9�`V����ݣy���~j�>j@ S皔����e����N�B��R�s �If�ζ�+:)�%8[w4�������k�z�(�㊚͡��[�z|�)m0��3�<'xu�@G�S��G�2Y��o#�o&�`�&0�v8�ΰ�3m[�۳,<�pCr�y�vM�������
���VV����%��aiɧ-��L�b�>�q�_�A �� qF�b�|D] |�fV.MkF���	(�kW�
�
{�|�c���2*+Ӿ3����"$�)��q,�{@�qnϠ�!}��i��
���P# f�/	i긑ZHޣ������&�����cƯ��d�p����w'qa�,�E	�u�,F,�����i�
����tx�4�P��Ky�?o�x0y����iQ\�Q!ү��CL�Ó�ӟbN[���{�'�m�д7�����ԅ��)���bcJ�gvnm�o�"+Ԅ3��{�+��Ӯ��]M�Ʉ�:&����{�	����ɇ@)#��?ć2��j��'����w�EH� ��:�HYȅ�.G�mN$�%��'eX�{1��٥s�\C�~��l��_2\P�P�z�x �xu�a�XD�\C�=V�� �T�347g���G�m��)|�iy�OC��
И��E�/CG�0���a�ηc"������xq>1@�="P�/\�c>�_Bׯ�?��u�� �G>/�򏪵�~�r���s�)¾A��)�y5���)���9��o��/��s_9)6U	��^93{\��:=����ڽ�C��q�ц�\��Q����TЮ/��ђ-4P��x��,�}mq0�0L),�e��u]�h�] dO=?A�2�k�"����װ�����>�D9�b��"c�Z�,���k��:�+�#z[�p�2.�*��{u��t�J���ȓ���3�WN�����nf�}xA���D~5���}��fe�@���ʗ��:ziÎ��{	8� 9A�/FR�S}�1*�'�JX���;C�%}Ň=�ɱ��*L_�fs�N\��s�HRv�L_p %A?jsv;k�xfYPA����~��jRn�ꡠ�s��<�,\�71S�H�T�
���V�L�@x�{c��ֳ����S �@[<Z"� ����p㼁�g.H7��,�����A���ňn�-^
�ãq�]���
q��w#P�ޱ��:�Ǣrhcڧ����R���1.ؼ�]ٍ+�8�`0�	�����*�}!Z83����|�U��( W���QG��%��f*EG�a�%�G�F46>]珋�g�Ml�綹���)Ɠ:�7����hj���u��NU���h1v�T6���h�
�@�{o�q��[�|��<�ݓ�T����a>[���x����.��DA�݉ޮ��%�����[(T�
�	��JF�䲂@4eT��Lb��q��hXO�}z�χz��Y�'�M��Z�t�Tn*���r1"�;���=.�Ǆ����ճ�v�$�Z6��v��ԾCL�'a��X�J��#�+��ͮ�����7���t��+��D����U�9)u0��)��V �W���������O|���h�y�;�ˆ�D��7;G9�W� ��x�@z{M7���^K���	Y2-��uT��>5Q!@aO�Q_�W���PR���_.��� ,�8����}�~3�G-�����<t<e�*��UU��&�x��s|��Ǹ�z˓P�7�{c
��$�?�Qy�t���Љ�d����̱�ןo���Xw�p�:��[`.ߖ��[�
���n%J���x��/TG���d
�����ӣ�V�T�1��^:~���Wye��>}�L��cL���O�z�T�I����6�Nۍ[M�;�\��<4���u�J���>X���z����V�,G��)�A��*�h�H������MH���!M\8Z�C�FL>�ϐK$ez���	au*�k�8F�ڐ�p(�:��`��8����Ax�'�������_Jڬ/���/$�3��