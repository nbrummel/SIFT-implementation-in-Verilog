XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��zB��A�+\�$���� 0�E�~n�
�v�Lz��0D��U�C�`u1�i6>�(��f6��A������Y"��ed_emp�J&�.�'ɋ.�S�n2%��x��`j�{$*�\�.yX�V�j�<K(U�of� =V�:O�B�hmU��LG7�g�]"2~J�瞁���U�<���+�4������*L�_xwھŲ��Ĕ��k9c�B��f<��b)�g|�)�D��#oCy���Z��r�$�˰�s��;���~SVH��7Eln�\$"��ni�i��2"�%�P�\z>
�%fN��Ea$p<DaHx��o_㸪G;�BM�a�1����险v��r(�P�����$��&S�>��J��)�&�]͞��������մgqὼ���� %�b��)mE��������}o�8�l�\�2���&j���:�ն�H����G��+÷�lߊڶe��a!�3�y�ձ��i��k��Bv�MJA�'6��W�)����^�A��N���}�>�����i>��cpyw&"�#�%�Jh�B��.��J��>^���F�x�B���b=�Du�P��U��`Uٞ��q���(��Z��(/`pk����8��.@�0�^�wH�@�h�㦦2����o�I�
��Z���zѝV��珗2l�'FJ<�7V{����Ǳ��t��HX�9��Ŷ��v���R��,L�#>���
%Z��|�iQ6WK�<����T*�hC/��A����.ZW�֒�9XlxVHYEB    5694    1290�xBr���\���vh�(�M���1k�RZ��$�� ��j��}H��N��gW�Nfȶ�0؈(-:|�n%l�BG?P{�t)S��E''��w�V!Y�h��Yϓ���ϻ���=�R�H��n�(�����"�6Qr�3 ��
D�Z	��F��PӴh���ͻ���[�[�	hs:���-��t)����U\��\/*���K�v��ĺ��N����p����m�s\���,����v캁r�v�*��JZ��/*��i��s"^[�}�#5)���X](��2.�k"�p��(CХM�!����P��/5\u�5{M�믰�d.�x��0x;��S#�EF���-{7e5�U�f�Ŗ�y~��+�t�i�3w��+R^M`l���*ݝz����K���H$uh���{�a�H�ȴ�:��>2$��"�>]�X+Ǵh�=�,��������՜_��ş!���Ї��ftW����aY�_���"�UN�[�b��M������*�*�j�]r*ܝ��&����K:~���7���H����W��u�Yϓ.2^�-.�����G���&�]�u!���ľ��U���;jJ��sV�Y�*wJ�Brt���n%:�&�P�#����j�������|�v�����q�A x�6�h2�+�?��
:�)��]�T"L�_DiG2��t<}.^�� E?V��j� �98������=�T�v�fhJ��E��g>js+��Q+�lq$-�h��2)��9'ƈ7F�� �X�a�.��S�s�ˣh��������Q~�\�\��<CnT���A{�S���jy_�R3�F�O��|g�v��,t�#'���f�ӷ��q�7v=AD61
V�Z� g�'	l!�	1� ?�،��(h���>dz|Zo�x���cN�8��B����i��Pn���
�ˤ�#��1n����w�N��1M��v��Ǻ�1�)y�)X��H9�!�V�� ��з
��]ְqG�U�Qn��	�L�wP�Z1v���B?R����Lݶ��)*�v"�)�Xn�Ӯ׃h>�%t7@���cbT�j7?��ER��O��`�dໍ΀!w! wUt[��eQN)i6�W���/�h՘5�,��Q�݆�s�$p%�!���,��hG���lʼ]�z�"�֔�)�\7D���DY�S�[��6��?I���E�=��U�A�Hɽ�Zb��0��Q*�k�l�+)��,�@��	I0_{5S�]�8#]S[���1pȾ�'�c�~$�K�����>֌��!\����,�:�d�����7|ֆ�	�Y�X:����>���:���M%![J��T�X��
�ۻ=�P����."�.Y�$��(Ac����	�� �c̗��Q�#Tp�o2$݄�u����b:ө�)����"��r��G;Y��%{dY+��5��G�~��2{��Z@) oq�s��t!�M������w "H��_���\r�z������9R�Y�B�ugR.(�2a�/���s�Ԑ�OQ��`c�&s]�m��y�T�q!�����sZ�1�M|�YNtBz�$ �[紻g.$&?��#V����`JI��U�iˉ,�k�Jsn�D)��0Pၱ�>�8�|���I��~����u�D>��J˘�J�m�M�>�4��6F~L.GP����/�ǈ�#���ڝ�$��c5�$S>;~��v��y��[��w�{�
P.tLrw���m%����%H��V�Jh%��L�؋�o3�~`bT��e�>F�-��P��7�2�M�L�/�չ��4�.0	PL|��&�N��7�T\��
{g8�tHߧ+$E}]6)tIEa@U*,����)��� ,j=S%���<	�*Kdx5�@�N���Zܪ/�+g#=7�<�P:T@D�jn�
�e_�h��L�4E ��ܟm�=���Ѹ�`�O�½��<X2d]�����}<�Zn� OǸn�k�2GfV¨��<�ξ��<�mc����s
���,[;�iI���р���v!̏��(\GW��n��h(2�h���"0��.�ʌ0��C"6B{pޭ�Ao6��u���A!09�kz�� ���6nOQ>/��V&���M�"C,3)��􉬿����%`�G_��0��3贽�Ƞ�X?��?�.Ԃ��	�v��+����
���f3)�;�V%�j]�$��bI�V�1 �E��f�`��ݎ��%�<����+�T'ܱO�7�u<������=rh�v�y���W�L������Ψ�� ��&���M3*h6��hu�Y������6��>��������QM��x�|3H����uحA���ʒ�(�4u��>��*��j����|�3!CF'J�'Ɨ�G�[~ ~��Z���[Y���#�����V�E�m�=���q]�OgV��*�z�&ؤ��Il����·vm̖:G��X��gc��I.Ņ'�?�}�����Do�3�����1���z�6����8��;���\7����_�~�*�Ns���O�7�E��:�b
��LY���U�J+9�:�Ux�?��4����s��h���Zj���+����RfG[�M,��?1�� }��M�D|1*�3�g��p&�~��|�7~F�(��4��,y��"Iqg-"2�\3_���3sT2�cB�ډ�:z��""ư ��ɚq��Ε�漛�<�QiDb>�7��yM������Ķz�����<�0t�)�$�Q�
��9�����fQ���/ɗ��[ȵ!֬N(!�:t'3u��M~��1l�pP��%k�;��l�{؊L���KxM��4��9���q�l	�L֐tٍ���A_���(ygQ�����w���9.9�C@�I9j�5o�Mg�];���}���v������Ұ >}°IW�\p�
JcR�F�K~[s٨j�|�u'�:ė�WN����U�'�Z�P�v�O[֓�eK��Mh�n*�k�i�ǿ=ТH��HZxZ���Xl�Ϩ�͌�Z�5�$6���n����F=4g�	\��K�ʾ_�U�83���Ze*�cy�ӼǿVQ;uҬ�- �0өME���%�đ�uJ���x3�>R�����6`�ά��;m2��qq�Pڽ�Pj���i�Q����/G1U9���,��ռ�5q���S�������W=0����a�nD�|�����ߊ��< zA�?ݸTn1����wt�5pM(I���C�ˁy�k1߹��\.�� 
��m$D���m*���U�7�Aa�i $�~�7���7����^��f)C?�M£#$� O8f���8��h�S����T�$��гg�o�yDXs㱪��G�Ln\�ud�I�ҕ-�b��7X���z��#���J���'�ujY��D~̇�&MT�ջ1��n�?�\�����X����s `w��.T�NX�@��F��T`��RD�O\L�4���˟j��ڑlzD�lV���W���o���к�����,��k�$!��՗$*߈e�W+��*>c�@��ș�gv`�#�q�#,�ǎ����ۘ�>��P�g��>�Z�ⓔDS�c��.��u����
�����Gح�P�6�_�&�ͧl���L4̋&&$\\x�o����2�/D-h�V�=�s9b���6'�+|ҁO]�ͧO~��� m�ҭ�P�A��R֢���7?��N��ª}<�Q$�.� b�ʭ�4a�Z�[<�̵��F!���5b2���� �ܙ��/�_�|�;��~�\v�P7@~8���~W��u��z�����/�T/
�ȇBBI�ĀQ�33Q��ꦁ`�!.�S��m��J��9|�P���{�A0\,��H̆�����d�q�H�#��U2�^��)�p��'��h���s0w�Yl ��R�AN�kn��
t�-�������v�+���7������>C��A�(b%.�[�Xjj�����s��~D�m	��� 2j)�Oh����l*���i8��ƒ��=�P��DyQ�O��T/;x��GaҕDRW��*���;"0Gϫ���Ų��oF�Z��sd�����6)k�4��C闱�%�4�RJJN ���^-9��zS�T^�%� X�����I��d���d�z��i��`8��d$&�F ��&�>Y^!`\�N�]�1���{�ʫ�s�Xȫq2��+�	�T�
�!;��0[nR�?�:�x�C�|ܨ���0N��_�2C�J s��Y`�肣~9[F2�=��%q������9�9�z�}c8؈P�Rc
J�[/��m$A��*�iZ�p��k}I��轶)'�$W˭g����T-�rO������V[#�C��*��*5��j4�Ҹ�[B�<G�taG�	|��ee���ŭ?&��}�B�M6�j'�P�9�х��F�ӷ���#��NI��L���7��6��X�������l�k�F�K����O/ɋ(ǋ�jz#
U|�s���t�К���f�Y~���K.-�`��)��}&w�PV"'[ώ��	�i��X��v�z���%�)�em �I@:��M�`	H��r=T[���>�Ő�kl�?n��:"�_�ݩ$�en�|��ri�y�,�~��|%ç�E#l�+�"���`\
�Rae�c;x��"�����U��/i�νi��1�<E������l�Q��bk���l R�ȡ�Y