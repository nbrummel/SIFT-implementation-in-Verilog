XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����F�\ 4`p�!X;kx���p��|#P}�p����G�ٷG�8��� @���'@�,c�I��Tqle ����}�=v>�e���?��e�<�����;D��y��`�"VX�����̿SLl�ށT����[�����+��Ƴ��w��2�F��@D���'��T*��rc��<��12�F�ʐy!!p��ݘ%Yf���US���S�ԊvE(UB��ů��bLK��eڰ�3�h"�﷠�tЃ�rG@���؃���CĻ�	��/CÏ=�Twɉ�
Um��;A�,`�}��=e�c��	}�i��M��	]����rj�C��$�[��4��.�=0y�M�\"��گ����~�Yן��vcb��ujN�P��b�����@%>-�u�:2��oٛX>򝯶=���+�~��	�HXor�μE�&��������b�<}�% ޔ| �����K��]�G�-9�ک�¯5�q9iPS����O�014�����a�fd�A�W�����B�0�DB�q���O�1�"/�ߣ��e��ٶ.��P9Iu5�#@V����ӂ���&?]�ڍ�#
��Ll8Z��R�6�6ԡ������q�Ĺ�ge��^X������!J�\���Sa�S"�\�"6.�=�à�b#����J��#Y ,��!mx��JgS.�p�6�z�\LC��;P���C�`D�l[V#�h1�WwUi��4���5�S@��MfɄ���L�Ul:-�-�AXlxVHYEB    4a8c     ee0�H�L�i�7���/��-�"�:A}�������}���6������������Ջ�K�0R/��R���|PEks�b���ݑ́�㚔������aZ�\W�Z�\iY�&!}�&�dpyv+���5���e�*��R�m�	7�ӖO��0�jj�0�v���t͙=%����z�M�iF�-l����3���!Cn!+g�k�'0Ry��dJ�a���s�R2�9� x��5�M&�PG�~זX;�u�U<�#׻�@?^V��>Yr���q��'z�y� ,���\o	�u4�^�E���Wz�E�����~B����P�k���Vзl&C�$ZECU)�	r�h��t!�GT�0�
�toT��qH"#@�t������6zua*��m`�J��y��(]t_����f��U�F(����-d��	�4��o��e?QB�Ǿ��]���u�~�F pz�g�e>�Q,��$����?�Bz�Xg
yj�;��p�;�t�Z�����~X�"~!�
o��:�Gg����Qc`"2=�����Y@U�A���W9~+�$��sq�g$?2��v�u��6C���[r��>��憕����E�|(�T��]B0,U�B�=����_X������W�JS�2��t�~o��ۉ�qח��G�?8x�B���L���?8௞�F&��� 8��C�&^�$��K|�璗Bf<��9<e �m�}���L�TT?�G/�Z��A���x�*��^^���Fz?�[);Z��1S1O��M�F�W�N1	hf#���@�Ңf;+U���^�Z����畒�X�����un���$�#F6G�iS��X�_�W1��@�C��[Ȍ�^a G\���i�%��Vٌ�p�Lv ����:�JުC	,L���I��ip�0`E5}=~Aʔ�&��cD)!���i���WF����z��� �(UܹU0�/�+�-F��U=��ӝA@���f%�|Nͨ=��]�$�e�4�2@,�Z5������/o�q�U"�o䐽�����E�\�$�r��fӷ���"3���'F�v'� ��lvo새��h�����>� um���������,�݁~�>�7O9��r�(+=<��7���i���ClBs������x-��5.k$�ϊpX�����R�͏��\��b9Y���*f��(jt!� z���/�Ա������6%�J��j��5Ŕ����z�o�=A�P]`z ��E/����s�m{�5��w�X�����}u��HާEQ���Q�c>p:&�=d��0��I�cؔ��9�����3R��I/��z����(�:N,�r�U�(�ƁQ�M�IY�c
����!���j�����W[�Q'�RB�I�z:ͣ�������*+c��*Z��������IIU:��z�TB��ug��T��(�|p��{����"�����WC���i��t��	k)b�'����9�k��K�Z�	A'�"�R(^����x�$z�!�s�\��i#���W/,\_9�ZvĆ/:��t��=�P�iY7�jX=s�����CWp�ر�E~���'B Ԓ���-��
W[�Lˆ��S�b�^��L������ٮ
*U����J�9p��>�Cv�6;>�m0&��^. YV5¬1k0㛮��J��zgB&&�,�(܆�]��Wj�Dȗ��DS^�t���M��'w���|�;I��k���������t��SB�������l�p��'˶����y�ۧ#���/�������6�S��^ܤ�E���$�>Eб�!�`&��:ᾌ�'�Q��QL���ܪ1.ҐT�A����N[�ec�X���e�"�x��G�}� bQQ^��i���E�@b��T�[p���{媺�Z-k+ixJ��ě[�v��\�MKg #i���蜮�����iSb��%O�?���'��5b�����i�	�qr���:N�T'5��M5"~[)�Z0f�3r@��wiM�pt��D	�!A`^ղ�rér�C*G��`�P�ĵ���Z�����ʤAֺ�hωX'�����e^�%�(���X�w�C��7pE��"�x ��=����P�s�q�1�U��w�|Nw5j"3[L ���/3& >�)�~�����}��^�>��Nn��
�l���2�q���4�(��|v������(���]�W�bm��L;}X�n�R�fX�<��"���G����#�t!ơ+c	qe��a����R Yl_<����V���D�����#���N�l����~>�*p���_���N�����6MG(P8��<�gU<�򞆆� v9��w�R�o��N�c)V��K�����s�}y��+��=��!���y�����VyV��X����a��j/T�U��i9�'2�\�e2�/7�~�s��%ؘ��
������*64C���%,C/�Dt���4���l�����d:������
|�a_2Pq ���ߖ�(8��1[�N���(�3c	퐏)�����}��`�l&�s�qљ4Ja��99}�p��4H	���L1��e���d�5�~d9�:�.�;봪#�� T�GO!�Vg*#yu-͞V�8�]��T�d��x��5����]�+����;[+�ծ򯃹d�lc�~�z�f,�����:sr��]L��.���] lh�8u�#tT�_+Y����\$�<|m�J)���.^�P���Vwsщ�!�����I�X24X��umal	Zk(����%ʞ��VfS��.��������tM� ���ou4�> ��g�X:}})!��=�\^ �5�IDR���~)C����RW�|ju OF��d���v��2�b�QM��FDf�fz�KSpt=��P��C��Nذg�C���`h1�տ�p�y�ǧ��*K�d/}Qu�_\�M���q�FLI���M9ٱ�.+Ô�a�7e��-|x.��s�׻<��^]����rWM�>)fT�K믌d������)�JS̩�d�Jq���4���Vk)�]���R��~v�?���O��<3�Ɔ��b,;M�R�(}�l�g�5�åKze��o��f�_!>$�4g�K�?-���J��������o����3ek�y��#��Q��4�_����8��h׶
M�AV����,ݭM.^�t��r��.Xt� \N���WU|�H��!؃Unǋ}��{!v�H>�M�qmp��R���	��5��ֹ�?�L��!ث�x��(��́Q����K쵔�/��I�J��U%G#lcSh��/��g=T��^�3&� #��{�a% Y��4����םkn�߭+sх#�˹b�KHUM�I�/�ځ�?�0��:O�?�]%?��wZ1�����g�O��=	�ZkcQ�-h/�[DP|�̵@QD&�͂_j��b���=ԘFT�Q�-�xmö��C��&��;N��5˶N5���_iV�R�/(e�U=�p0������ﰣ��6��P��,Fv3Nf�5����4
5����7�;	�5k�Aok@�
�i���P#/
�_�p[��8���O ;5�4�{+�XjdQÔ�����U<�=anb~&X�9)��/%�}6�/�����b�L�0�����{�Φ�ID�΋PDȔl,K��24���8��}��-���A/ƅ�㛹�nʐU��ž�IhzI�W"2����7�:7�Ȓ"�~�G��;� L(��jw\��