XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���E7���ڑ��������s*�'-O=���#Tjg�nG������e��{M����Vj����t6�.��Y�h���Q S��/��{�T�*~�~sҊ$�b��'�x����Z��-du�r�yۇ��G}蜬@��ޖb�@���%#����)}�Ψ��͸!M�	�'E�	�O��/M~�̣�v���^}�{<�ec��F�����矑јUE$���ٛ~��;��s�u0���3�����)���h"l O��;�3>�A�s%���7/�ͮ�i5mǚ��a*vP`�:��>2�^l���,�q��٤�[�0p�0X㙷 ��CL��:��������j��$"��?��VYL}�bg]d�0t3���!՚v<����+3�/H�4��+pt�a�D��0�t���ؠj�oj:�v�X��z�"�������Eus3���ɕX ���>0��s�;�Fi��=!
r��bt��I�q�@	w+`*Z螰F���e*i�ia�a䣑g�D�S�.{V��NCSj�/��E�`I�i�Y��s��5�-W�H��6���Sq�	��R���tL��s�B.A,G�����V�A�����'g��ݫk"Bt�	x�SH�b��@�B�q������Q{��-_^i�����V* �h&��ڿx���:�mߣ5��[r'�I2�����d�N3Q�:�2�&fs��w��2�3&m��nf�)b���7��1h�d��dbi�@��؟)�XlxVHYEB    fa00    2910�Vp�����%�2dG�G�Y��W{p�D!�ƹrQ�x���A%:��4�/�%'�<�����0D�SV.|r�y��}^���������8�q�o�6�3R��Ӗ!� ��-�8KX�:��(8%�'�1V\��
!:B�ǳ����i�.w�h[��Jk��/�'V�{��"�cZ��/�˹���!w�&~�9F�ի�z]�)��i�tS�Zy�{|�e�1��@MU�>��vD��k@힝~i�P���>N�Ķ �6��ݡ����59H���c/���}�J�:����J3e�;y����ب ��LexE���i9vkĈ�;�;�:}8�O�p*4��h�}���s��W��'Y��
=;�F�	�6���D��b���̔L���� KF ��=9v��~�c���$��5
�?�ͷ#8�V�W*i&�:;���[��ܗ8 K�@�/���z�`�;��A��7�A���㦅�?#(Q�%���C�H�%�x�.I��.�N�Y�z���l�b�t=D�a;f��N�U�`Ү��>SC��]��X��r,��͔�p�i��*`�ڕys���鈐M�=�%����k� EQ�08(���?~���|�Hn�D-���l鋉��btW�T��@�#�c��3�Y�{c�^ø��jk��ӽ��៰X��� �;5$^���{���4�������n�X^�S�<aè�X�8�F��6=�5Ϳ��ŘC֮� �`u�/���/�<a6y��m�-�����[;As�.�lF�ǧ�uuwRΤ1��S�B�����ΤZ�׽���d >��h��-�oM[�=n�L?#I�!$�W�k2)Һ+Ws|:�^@�ha�K'z���$)IG�M��cNA�掽x͚�q4� >c0�J2"�Y���=��T>��Z)8�� �n�G��c�/�Uچ0(�A����R��p[�'�hY�:��s��W"��`���	2��a�V�vW,�!���ʃ��M6VV��T�����hR�}7|��BMZl�Z��<��g�r��-@p��4/u�N���ќ�d�٘'Å�h��P�����(@\v�[��z5jB$Ř�$�g;�t�0Ͻ׫V����������I$��pR��-�z�0�rlH� ����,9�0hR�=����h��`�J�F�����Dz��ǘ�l ;@�P9��^�F-|�j�/p�=G?i�au�	4.�h���$�a��a<���slw �@;?���V���@nH�]!���F�|��*):������a�4/��x��3���w�z�+� 5��k�ك����B�7A3�ῒ���*^^?ձo\����r��f�u	��Y&���*�*�k���>-�2+��lmNHF����|(��o���>_⃕�,Â�9�V��'4#�W�m=�7�#5��>k7d��R�y�(�[0r}��z����G���w�R�'�N��j��RO�&���pX0FQ�uk�7����c8 geK�� ���1Sb}�ι$��џ{��\�\L��՘�+z*��9��'���Q�i�ft}Wyy�>�ui�qi���g+���*��G����ːI����i)��\e�f]a�)��w�)G�^<tp��Fv}Y�{�O���B9�K~�w�,,�@�>6����)�6��a�,�é!%|�%����D�~,_�h����ϣ�\¦�1A��ט�g{���{Y��ʗ��3���zb!^�7*@��	� &��/�Lbl�������S��S�����	�*zh���r\�1{��2(.d�|�!�y�N����§��fAb�4M`S`��(W�3����G�B�*L<�8���Y����)�(�t���@1�7	��).���h~DRa�ڽ�`|��l���>��x(@��w�B���M�m=n8����w���t����	�B�|f�`w��w'�&z
�5�
P��҄�7q�ft��r=H���r��+f��:[����KP�H���dW�.[�Ϳl���Yⴐn�W)�}����@��:1��~9�c0V��'��/�kכQ
-[��j=�O-~/�o'P�D9��(j���=�B�WDw�佊#�TZU��,��2w$�ߐ���S�H���E�~ ���~�Z��E
-�nl�9��|A�A�Y�C��/�������04���m�uT�m^�c�&s�G�%.��7QBy'�.ڶx��h���ٽ�iy��wT�=��3l��� įʴ���X��5	�?.�]#>�����D7U^��͏�����Zx��Sg��R2q�7�01�����U�=�H*WD�H�.��="&g{FH-�߫E�_�4����mRxF����.
��"��Fp~����?�e6�����K�yoP�B��pִ=��稌v5��q��[��{��xY���/:@��8�z>��5��0���MP�Y6�_��!jx$'���� 'e��n�M�$��qߧHH�}ti���~�'w�@��zMp��M���F�U���jۣ�z���5tpzi��$��倥�;߯xi2����,=�,4,���ٛ��_j�c�л ְV�fc���]>:=�ӚǶ r_�_�&HFn�m�,�0���p9�P�K��و�v;���n4dPn��;��4t����K~��4F�:�����㹥gK����<����vH�w����D��!7������k�V���I�̩���Hy�8L�ؤ1�f�C"Y�TD4�z�ф�)z���i�J�X�_X����aD��<+�p-)�lM�=���� +q��޺{j�4���3�y$�	��p̴���ϙ>�1:2j��i[c;�6�_;�Ɗ��$�C��G���T2w'9<��G�=ʽ^��L @F'���[�MZ>���^��4L_�i��`yF/����L����+Q ���Ѳ���㍗Q,���u�&#��{�MO.y׺�!@R�ux���7�=���glE1���	*����w��դp�?`��=�� �$kP��Y���z����y?�o�~��;Q $����S.7^n���F������)c�kR��ӈ˃(8qqg���fuw�v��7Ju�J�;gK���@���R�V�5�����E�O�=�t�MV�M�ʵW��EZ�4,\����ĸ6���G��L�1�c��Ü�f
�� �P9�S|�3��q~ޞ¸�'�� �wӪp���Vވ�>GL�T�,$�ݻP1E���l���*�y]��xj+=,���?B~��"#���w��&�1)��a����P:����\�|�7��2=�,�V6�>uU�Ձ���8Qפ��_�_B�\�Z�'��VA�0e�����p(� �ؤg��/�z�Կ��1�����V�Js���F+�ʑ
�Vįm%@�XÆ�i���Cl��b��ogE7�����f5_)�?�	��K�Z�	z�>TW��%�Ց`v���>�"�R,8�P<�k4�t�%,e���i��M ;��2+o�\��.��9v��%}j���԰��qqK��[��ɨ�m�P �-����W>���� ��bfЌ�!l��x��3A�g�k��I�2�5\�Qz ���Fa�`1�F������d���C����>w�F�77t��JgR�<�����olA��ƞ�z�2�`�V}��E��<Emj(�C��t�cr+Q����"���3��%���%Trڍ��aB@�@�n���=�[#�<w����ZAޓ|�w�ߗ��W�3~��A�+1H<��h
�\�̠�-�˗zx�ꊂXZ��s���Kv�m-�$r���.O1G�ٞ>����k�]���ߌ�c��Y�}-����ԛr��@`����E$����w`M�-���'��/Q�U#|~�S���,v%�ߛ�}���1��	�"���$i�zaX����M\�$3P�`G�����U 0-oj~'�4��|+�i���z�� ���ecIf��q���^G��n%���x�a ��u%��_h�7��Y1;g�O&�V��ip�
7�V9�{�פ��⒳�Q����6)���������b��hK�0�3�
�g`��&ݩ@XNm ��|�#T@D��w�*U�~��K�Þ���TO�5����Z�%w�:؀�9
l��GV��[<H>�����.��ۜ��u�M�`��ﴊ,'��N�-w%CC�=[�������UqT�=sec�@Ԃm�?� �Q:.��l���L�Kp��w��-A�T���,:j �|{����I�P�Y~�4�7ׄ0�y�e�0�rIM��4K��"�B�G3m���oN��R��sZca4tu=��������J0pov��/Z�J%ۊe6~Q��z;��!�jKO@�ˬ��;�1�J�>�RX9���kL2� ǯ�,z��ӌ����(_Z�}�k�-�����|�5h�H&+c�G���b��ħ���/�xR��H+���.5���S��"_���r�DI)�F�Ɉ��ط�6�G�������ubb�R}����niP�U2�G(DY��]q�,�]k�P�N�w�q^� �m��]I�p]��i�T�3R��u��P7]ϓ�ލ��.O������,��ʝ_i������|��4-��2|�ְ�2���쫑
J�4��*����L�����I
j����ku��Cm֛S`1��,T30@�=ߒ���HV��&XJ�rJ�����c�ZV��H�Y��z��:��޷c�o?|3q'X".��<
?�������#�G�	�\E�hUU�i^��ʈk9��,s��n37(��;y�Jv	j>���F�|���e�z0��Js�h�������y���-X����:�E��Ϭ�mg��މ�1d�G#u�*NZQ��ٜ�
ĳ����W[�S7�y������2_E6��n}>�A�KK�eD ʢ=>�ܒ�滅�uGc#�Kˇ����EH�m�v>����̻��C��/��Ű����������Ӫ;�v���%���/�ݱQ֝��Q�a�[�������~d�����J�����(�D�C�_��̷uL�0Y���ߩ������٫<�Am�U������r�koL����vZ�Ǵd|B��rL6R�T���d��)��`�=ĈAsm���n��::£�'����2c��{l�s�s�����#�o����F�gi�V_� }ᓫ!SЕ��>��{������z�C�2�vLHE��n����,�����f����W��%����r���0�{�I�h)��a�V�ӿ���OY]
.׶��C��k����PJ�7Ee�a=��)1�PD���H���!"�t"�_�Z>�|"ԺEDatl�r$�L�w����Ώɋ��v�h��c��E6(G��E�U��O�� �3���3���l>�8E��A���2K5Ƴ�Q�9f�-	ö�����6��������A
@���������?�Ga_>諄�f�����#:���"4���Z=�%ß���Dt�,9Wn��x�����&O�[W��FR���Y���ʴ�T���Ǣ��R�'�[�T��Ky��6�w��s�i�O�RR���)��Bv���<�bj�<�G>⁷�s-c�浛�n��� W��R&&��MXy�iM5�O6X"�x���=w��P���6S�l J�M�s	���Ue�Q3m�W��p{m�@�.��n���ř���~'���@W�Ե�r��C�TT�����Qi6�m<���dl�����I�ݽ�8f�c��\�]��k��QP�_�i1*AH��m5�7��K"j��U�`a �&k�ib�� ^�3_������w�=f�҄֊��n|J�a@ _�?2��7W3��XzD�1+A��pߌ�y%���3��_I#+�[��RF���k��C�u7�F �f�2�̄A3��"��R�⒰jD���)����{��z_�CטڅG&�`4��%�%��,��]O��p�|�u�V b���^7�[�ܡ.���
I�<���쬚i��@��R�1/���t��T�~���P�@���C*ÖAFב~��&����2�k��䵓��Rt���,̪��#B���>��˱a  ��%I�F=�#eb;�y�Ǝ���88���m;�jw��q�>�����[O!�~�3Qc�����o�$+���<��cq�Qnd�9����p�/���9�tΑ�x��'��a�<74���ʭ
�E�|�ԣZ��L�/j1�(��v�U��{����l�R�h��
�yQB;�����n�����'G��x�vO�f$���}b�����7>�CI�Z��l3&'i1c_Ө��'nH�-K(�x��NK�ښ�1��E2�Fc��q�O���	Nfh#�#�As#@�).E�vf_��������e�U\޳0�z(�PF !����K&wZy����a����E�E�8��P4;��5ؒ lo��݄��>���ry#!\�1������K�l�bt3�ք�
���U�F�B�=�T���ӽ��v��_[���[�"�~�v`�=ӽ�C�2n}~�� ������y�К��Z�c�7��GCߖ>�b�$g�m��DQ:fv�v���S�Pۻ�qaf��ӆrΣ�-��Sh��\���8�B�����+-P��M�
~G�h�q�Y��sZ�K���Td�0�������Ɏ�<��������π�~d\�1��`b����9�<��i�tAz��Z5r�x�؜��u�}����bf|�<��^�>W�OyJ���RD��U���r��X����}�!e=\䦎����ۺ$�Y�]��
���,�w��9M��`,w�p����h���B�;�@~�=�J�.��=��W���Z(w�}k0���f^\��5/=y'M�8ā�>��[j�m3}�Y\����C:Z �4��@��4`԰"l{��s�kz��J�Bg,�}���EH<���eqĿiFXF���}g��oG7|W@��|���]��0�m��9O@� �����vmM��$
�>�1jW��_s�\Q���_�O����z��mɼ��gb\�44���t�n�
����C�r�
dĦ��G�e�D�-�u�&�~'|�3,9@WRk6�t�-Ozv�֫w ���j	��QV���Pơy�-,S��K����!w������s����zh{���k��,Eh�Iñ �<2ܶ�U��JY��!���'c��}��am��~���ר�qC�k1��_L�"Xf�Ѩ�Da-�w2��L��җ��EH<(V���w�5�����Z�8�G����%����iK;S&7g])<݀������~����w͎�h,��ވ|��Y	��&�Pu���p"LI�l���"b�q�^����.ۑ�����|��%����~�H
Ψ�-
	PS�Ɨǖi�%Y�&A"�b	��}����f�cC�fn#��nK�ػ�B|�%�(� I#l�_�C��h�*gf�~�N��A�3�5�X���Ą�k$�.����`��P;8!���Ͻ�*⅜kJ�(ڡfY�eww���/�������R@��@��1�>��7~�
4�;1AB9��X�ۚ�{0��~�>�S�%��d��p����+�5���)1ݔ!Q����+ߢ�(�{.�g]w|u$~��em��C)>eGYm���gryw�����o-]���$*!�?4e�B�<yK.���hT��E=�mM��Y��	Y�P;4���t���Z�S��J=��.�<f��:�m�G\q�Fiԡ!S�mg3PAB�Ր�<[�/�K�S����E0`R�\���7'�S`�D��I�m�-�l���~��n�ܷ�c�[\��#yfNr�e#h	N��������_������0�ͯ\�a����n��`hq�lq�(+l3bF�ݸz%�gOYd�s�9�B�U�:1��fk�t��;��) �(�.2$?�� "��Ό�gzW%���-
�ƭ�9^8?�!�/T�ê�{���uE�����~��o�Nq���
�����w̴�m0�S�* ��Op3��zX��~���0��MLr͵nu�<��Nơń�B&�a���;4���ua�oVCd����`���|Y�	!�l���(>.�E^4�W2�|(K�������v�'`�����3���G&� &�x;P�Qo�#���c�t$E��\Xk��Va������t��pB��TĈ�J���dk`QP~�3��Ҟ�n֍�V/
tUI�hn�4�|�߰�:��<���{���A����`�a X;�UitL��+�C9B�W��݈ڇY�n�/]��H�qX���<�~c�o�[�6�<6�w2���Z��Q�j��?���ߣ����<���d	�D��������T����aoYׯbmפ�c!PbQ�ေ��;�ԡ!?e�Ƚ=�Elc��1A�Z�qQ%Rr������{B�8���c{�Hj���\e?��{�o;�caUv�ꙉ� �jZ���P���-료���T����Mz�Cz��e�k%ְe�H��<-�
5�woģ* h�J��۾1b�LG����RX����pf�����}���pєG��(�Ff�N/�3u�N�jg�����śl>��m��ѽ�'�]�^ݤ��+~iV��`ȧM��� X�|�^�/��|��w��BA����[Mco��as%[|��I�<M�<)/�/�����{�cT���G?�E�'ӑ��U�J��>+y�J|��iq��H&�_p��8:�d�Y�s�n���8]��!�^����P��f;7D.x?�i]|�BJ�[���	�N]2��be
[��4�7r!g���a�"S��d܏7aM���K�M�Y���0�/~Agy�.�Ao"am�$�&5>}{L��<&*���A-�ۻ��h�����������:I�"�Φ�ʊyqDMj��]+W�&�0�U�-���?:Q����{B(>����W�,Ln|�m��0u�� āi�e��rf���ن���R:�b�1�9�Y�w�D}�T7l�x�2/������K6z���J��|�h�U;�Cf�2�3Q�l��M��
&]�'oJ�����\��vÕ����K�\��'��Y���"��/0|�C�1�4�|�]`��I�{1��a<���c���B�AW�}�(��fp���^�#� :)�B�z�U�>&
��Yђ�X��n d�!�`�_N��C\���D��7ୈ�?�� �`:�j{�j��_h�/S��Q
�����Ra!+���/W~O�h]��%T���*��q1_ �H��I��E
Qg��nu��z�tC��R>eJ���k@X>-/A �p��F�0҅�A������k$Q�}�n�{�׌�Yw�8�XT�v���f�X8������cNpj���a�#��8GJ[�.�W�)׏�������O��mM�8�*tSA��Z,��'�����I��s]����Qv��	sÃp��&�?�^�,�F>ķ��9%
��˃��}�ĳ��2��~��>��QUo>ܐU ��!6�û�g6楄��L!���n��1��~^�����{t������ou?�Y��/���,��㯿���,#;����-D�������pH�%�#���J�-��@WF��B�I���!���t��j�б6!�ݫ�Fhۺ�cA�]-��� �|�;��]Ф�KQF1h�q�c��JDV�\�B����J�t�_4�P���i��o��)����jC>����Z�ݙA��~C�v!��9^�5���x��N�B`Xu�G��X�6�;u��X����3*�?���^���s$��	�NY"��WooO���hO��݁��{�an�£7A�V�F0^�Z^�/�6+B�ʲ.�V��� �3-e�5q��
��K����G��*����׈ۃ�gpN��P�[+�E?���FF�p����������e^+�dHT��D\�/���ub�K�mg�B�i�00>5��Z�#� "����L��`��ke���H>X�3l9Q��KW�o��[�(��U��|�D� ]��څ���?P�����؍�X�А}��!Xf���0&�j����y
��͛ϟeXf
��l�0��pq�y���H�=jMolPR��j9�ض.nwt�(Ug���E��EO;i��آv`4�m/uS�Į�+�B�r;۹��[��Z�"[������XT�R�0�x�ق�S�� J�*<٩� �=tLv,���;�5�h���PP�����5��kBx���u�ai��������8�)x �E�}JC&*0V)��P����^L�a���j#'�Gq�XCu{4t;�v��;�A�)#?�h�d5K���B�\|gJ�2F�{��IGxn�L�XlxVHYEB    fa00    1d80�,�M-��=��uo���<�z�ܕ�
A��U3� ���Sa�O%@=*)��s�� '��:�cx��)(���Z�)�#܂��ڋk2��]���l��0�t����C��	,��8��?
��˟k� _<��a�uc �C&�,ha�A?��EЙ��'/4t��Qu�9y^ZM1��I��ܰ�� c��֯S!.�0�2~u�-d���
6m&E�c�K�����~\��u63UP7~�,�⛃��x�ބn�0�C[��xP��z-���(&�9�}9^c�A���mQ�Ś���"�~b�B�oBYD��
���F�z�t�]!D����ə�)����y�K�\��j)�ӝ!��e�4Y9���U�n& �;c��\ƚ�x�F�C!ys�*�8���ux�z� �M@[qiWM��*�D}�P��b�JV�	�g���]K!<�w-<Ͽ���g'3��]$G���J٥����LC��{���V���=��-��e^��@��^P�~n��΅A�6�¹����9��h]�D`%��LN�~5+���䖬�%c�Գ�¯�_z�O]���D��xh�"s~ps�P~���r�@�I�9������jഠ�bIp����i��6��obt~�P�rMNW�|M!M�h�&$�,�땭W�Fv��ژҺ���+���r_�v.j����� l�[���܍��=�k�	b6dtIC���/K_X#��2 ��[��)E	��Sw�A�ɋa>{6O�Y�Į�dJ��R̕B:�磰�H3.L=�H`����~K��G� ��&��c�z�av��O��s%�4(���C�݋ ��� ��F���D��1�1���o��F�.����=@g���$��G��k"�҇u�[��[<~����m}���긞�A��p�p2졺��hD�L�F�B/��1Ұ���U���V�(��4<�u����4�y�;�/������A�����_N���T�|>i17��`��J��<V��ņ�3�@]U O<>f�Qz*�2+�a}�d��?���Y%�<�S�r
Ǆf�4-��S�x����BX�����w}���DpeLJ��+i�e��@R�d�q4zj�Ǳ��V��'��ޑ����*�n��|&ѸA��xot������=�
,P8� .>-�_>lw�}j�����z���k�J�R�pO^�V\�DW�^��*l�2�-�;�Z�3l�.T���t猺��|K��qաǳ�N���w�|��mQ�?Y���; ���g$9���M�0�؀�_��(������G��4����z�6�ΣS���ʄ
�쑺��Z��l�D����a��zA�P��� y�)���yn/���ǰ1�ю��b���@ h.��E#��!i�jz]��@B���g�!�y}5��q�=�2Sd	D��=p 4�g��t�C�i� �Do��n��n67�#Y�A��"���Av��(�ɘ����u^}�� ���ж4~�N����D��14�l�� 7nNE@/:�^'8 �eё��bE��+��m�lAp�J�S�;S��s��4��� g��>[�|����V=����шr�/�0g�۱i�o 㾤��կԬ"��4m�6��-qC�'
���cq��qP�O�|�Dz���K��'�iz�nn6�Yˤ�Tn:	FU�:�H��w���|���=����ҥ|d���lS���5��a�:1�RG��_TH���+7w�T�����������B<Rnr���h8�6����)�/��iۣ�8II��ۺ�wu��� �$�k���_�?��%i-_A��������(b�ۖ��a���=`� ��u<S��y�̈́�'fS��Gܸ	ؙ.�HX�x����L;�w��7�	Od�?�
� ��A����eZ^��T�I�|Mh'�t�J�R{�^~�������1�!r�	Xu��P�
��p�"g�]5�M�7<%pa�da�)�ᡩQ3�t���� �o|\+;M�X���(����� 	F����΁��F�괺y��k����c�κ��|�SFxlP��E͠����W�)�5�򑬏�7��Y��-:�K��*'k��?�=tT�cX�0�u����ȃ�`6f�&�G�s8g[�q�|GLOh ��F
ux�;%��5��$&������������4�mQ�wP���Ƴ����Ÿ��m������D𳢻;JhMldyO�,��'b���DЩ��j1�/�2
 ?�}�V��Wjy���L��j��o<b.��.L`�TJ77�^�j$lj�˔�YI�"��t ��taĺ}V6�,��)uĳ�GlBv�>�K��:ؗ����:i�(]�M0��������K��迓��xF�-��ps1�E`%n���ӎ�9h��t��`Fw4��~���4��ɏ2�,�V��< %cO��"�2hb�@`�S(){�J��ୈa7rD����b�W�d\��E�7b��6	�L^@�Q*���݅�ݟ2_{�-�K��S^G}�`Nk
�3�\UG��p�I\l�ːh�
Ե\L�</F`�]&�0��j�u�����d=X���#c�M�N���xd�R���z��qu0�i�@+���W?��&<���V�Ѷ����0l�!����e���ݎYa}b`d�ː$�s9o],18���l\�^�-7�e@,�9`1`�vjq�҂c(�����^к�5PF�L7d�m�RCv�R�	��0��\�ͽ�᠛甒qO᫿|�Re�g���(���W*���6M=X�^��n�,ST: $5��a�*�Ryp������ng7;,:�A���
���F�_�ɰ��1e�)���������g'�r(:��$f(����qg⩬V���;$A#��/;��l�9L�M���̃�К���:S��=[��L��\��Z�dν�:�����~2�!\�����7��-�D_R� �n���O˸��S�ۢ-��b"�W(;����tŃQ+s��+k�Ź� �q�M�âI|�甈OZ��͊K#:��1���q��#2#Ϊ�W�#R�6�d��7Cg��yUnn@�1�w��\�<S7~�UYx�����,��~E��%�yeCݏ��U�H�؍,��v;@���|$)�3��[�9Q��rb���OL�%�9S-�Q�!]~�b�W]�RAg�
&����l�ݗ�/�����Po�iCX̥
�_m)&!�(���BN�����|�7�ơ�� 4n���/r穙x7d/�K�Emr�i��:������_�����`O����xnE��i��l�)�Ɂ3�Z̙Ӥ��#�M�W��7��+D����uiʁs?�T��t��J|��M1���j��g�X��v��clE ���D<Q�z�*[�P��R��5������u�Q?3�)�o	�������������9�z�Cp��񓘐��E��x�[ɟ� �)ː���YPq�@��>���sXs�|�(l��L�gb�ދ5�PW�����z�8R�C�F�悠��Y��R���u��� J�c�����`\��#p�}y��Wu��b�Ak,�ez�/��z�~཭�Q�+�^M�kw�=kз�3�~�6�|=0�jf����� �L���P�:�?5��5�	C��	i�*���ߖ��|֡�|G��V�T��K�E}z��nU?�e��09�P4P'���ʂ�T�4� @e��6B�?h���H�����I6����
�P�^0���9>���yh#�*�Ы��O*�vH<�x����(>.�DG��Mud=,�sov�k���>� �1X�͘�9�lo<������#�V w_��s`%i����hx�L��'��j�8�pϘ!Ubo�k�4#y�����+��_�x(G�eB~��O2�'6���:�A�`mm��Ax�?.B�x����b�/�Y?��_Z�§Z���Ǐ�C~c��N�����ʏ�|I�$(��f�\�m^�jL�7�Ҙ�-��e~�����F-�E�=-�?�'Dۿ�)��|?�-�ƆΉ	(�I_�5��� �YE��UEf�Ϥ'T���=<��a�6���������{���bk�x3.��?K24�hɫV`E��)[4o�{����O�R�SJ瘔�ZD}�a	H��w �h7�Q�<B<3���;ۓ��;$O�Ǌ����7��/ir�)y	�ҟ������u�����E	C�#M�9���:۰���C�5=��0$���H6u�1���Ԕ5��� V��rO�`~#Tu[�����j4C�� n�V����X�tJ�Ӟ0�t�2���n"$ks�(�3�6�0x�i�w*�Z���#�P��tu�dSe��i��k�#餛�Qx�e��[cxQ#Й¨��3<�!-P��R�f��	vXQ�u�@n�v�lT@wN�IH� 	�~��P�.f��}��a ��� ��x��ɨ�������zL��-W|ˊӷ����1�ʿ�~@��f$���}n�C�~��M�#��C��-R���������PE(�6{z}O�J��`�q��_4&~��@��s���H~W�L���4��3Ǟ>K�1��K�^��e,����#ʉ��*�.do�!����K�x	$B�+_���2�ej���ߧ:�R40;�yr#u�+Vl�k��j�K��m?@�Эp�����@��.?y�ě#�{~G��uz��'�{ j�1��ى�A�7�DE�_Z��kR�h������A�{�
C�i�0ZEj�{"U�d�a'k�d�sj���5��x�K�:��e���N��,�V�
�e���Y�����"�H��ӆZ��ۊ�W�wt�q4y_:6�T�2#�Y��)VL	ֳٖd���u��l>��>�7=��D�L�[:nZRP�����m��T��D�IC�~�s;��=���w����?�������5-U�j�$Ix��$��T���1��z���Q1��3>�J4��Э�G�/˟�H}�8*�4�*�bDD��6�O��}J��Ʃ!�����T :G��F.�;"���`-x���.x����}���Cfv�%`���R���Jɒ)�^���SXLg� �X��];���ǶΩ_�𬉅S*;5�w�� %��b���f[����"Z���ux����zJ��s/�T��a���q��b� ��[?���N躸�`��:*�b�]��)D��U`���J�]A{2@��C�c,��K�+_���DVk���k��J�Xo���j�M�^J����3�}�ɞq��7	�e�i>�B�
����g����R�ko�NG�Vb�BÖz�F��!
uKֳio�wߦӶ>�ܶr-e���$����	���u��E{f�N|��8�|]aDz�Yq��~��k̝�N��g?D94PD�L��3v��G�}��1�+�7s�Q`���|���z��CL���	���r�B�a.�ЖH��M^���m�����5Є��o,��+���@nH�l_;�!W^泲�>�h�M��*��#���7��)L�sW�P|i�Ŋ}��s�:����K9��of�ֶ���
T��n����!W�+�ɂ���k@V��&�Z�l{�����u�m���_
���{Ӕ�Sk$��������B��aR3_+���3�R�A�%I�=`����L�Ow���<���5�7��.�L�����uI��Nu��
<P�	@Ė��#�_Ѝ��[�y�/�h'pcb�������wo;� ��[�5��$���GF����Q&To����
0O��d� ���/@��� �O?�j�i%��b���m��P��(І> )��u%հ��x1�>��̣�qx�P#ۼ�k�1��������)�bvY�����	�-�?w]�K�F�n��v���(n᪬"%B�jˌ�נ��_�ʱ��;[��$���0���_���Ϸy͋�Jx��i!J 2�#B�Z
�"��8X�e��d넍!��[�X��gRhE�_��WR�[Z���#�\*�Lнl!��\����ԇ�%��A]n��}hM�&��Y`���Tbf�͹iz��#&w� ۽�k�}|��3�t�����y��:���?��G��U����i���ƭ���f��j={�ޒP��j᥵�$Ғ�Ҷl������8���R2�L<��j|39� �8�>��8�HK��*M>�e閉���?�x=�D(���G��I��A��P��,��O���։�*�_*[��� �5�:ݱG�n;��n4�w7pv�i�ۂ7p|��tcL<O]�Ђ�� �Zp���Ǫ
�V��m.�)k��*(��<ݗ�;�u;����v��5F�8�l���v�Ee�O����EV��PBʌf$Y��u�uħI��Q��X���Tȝ'}^�7N�6��ꐸ>�:��&�.b��3����P�#O/�K��q�n�pT�����DcM��g�g)�š+$���=�y��|�������ȵO��&�����wA�b�	6dt:��̉�Z����K�K�~��K�U�����ʞB;�Ā���dP��E��~���[�5]tB`@R$�\��&�M"��n6#%=g��yr�,�ˆݸ�N@�n.�"�����5 v�%bK�6�����U��S�KW�'���y߁�w�5p�껂�o����6�$�����<F�����7�mյ��A�3��nXO��N.`�/̛q������g"�؉��5�H3f*}����Dj��3C���/����-⦨��us�d��  ���9В+����c�mz�5���s�2��8�7Qt:��M�md��I���+$N���3��"#��.��7�U\��>h,�?��ɟr9��Tz���0�*�W�V�P�dM�q�G��F{|I��a���t��:�/�~Q�Ց-���Qn�dT��*y엙u;9�=3O�H�0�����"zx������;�մǠ�=��;�� ������;��N�J.gF��I4S'��J�s:`k���k̍�,��>���P�@.`�o`*5�����K������y0C��vBa�b�޷�ݘ��=��m�C�����R�H��*g�"�'Jv$�񝷍t6��R�o dWNE��a��a|���[��e�0W�7�`�jz�w$碏�*�����7L�2�G6��E ��'4����݆vKP)���X�
�Z><٧��n���v�K�~��s��	�C�U�M�W_�th6���A>H\:��@��9�r�ё��hXų�/;��u�i�|,�m2 ��8�UYC.���*�*>=N鶃h�:����l}GZ�X23����(���
��km�:�u��.������i�4��L�+ރ�2𠣧��1[V~����M<�|��Z�}#�k�$��> �v�����T�?f�d�`*�R���XlxVHYEB    fa00    1dd0�-�jp�-S��WH�Z6	o�E��֥�]J�ڝ�K����ݏDј�[�q���������^��m	D��a�(�I��(� ��Kx�qu�;Lg��E���4��e�|�NU�C�����Ξ$̓w�`N+vw�5�$Q��}؋�ó�&��VWi]��K���)��G}w�99��<���C�S�����i~�a|T�u)Ӱ�T#����^����B���o�'�( �%a�6R�=���G23d���ՇU��cQ	Cc*��H� ��إQ4��7����@����h�7�Q��/Fz�t��x�&�K�N���G�7]l��ۛQv�"k���`eN����9^����œ��.u�����X{d�`��ѥ�5,���@לip�|��O�|G!��ec�׫[���/1��X�qj����$T4�؍5���W�O)��$Ƚ"���Y�9J5�m�|��Zո9<�q;-�$�/�w n���qDfKB��h�����'nN`D�<a��[�M�ak!�#�r��sx=)6t�� h������/����il��Bg)�YӜءEű�U��	��٫C��	���l�HL��D���aB�V �il�їϭ����l�OicϠ�7^���S'|���>��S24y�d-y� �O��K���Ǝ�8��s�$0D_�6�iCn�2�+���")�1�
�ENV��)������y�"��ufE���h&���6�;V;'��1N��'����Jf�a���(Ϳ<���I["}�Wmf�w�8��F��3%��#Baڅ����u<Na���9�ݘB��x����Jw
�5W+�
�!T�ӿm�I���z����xP@h�{t��&Z[�ęG=�';I|�tٽk����1 ؟ ?3C[�8������%	a��A��	��V�˱�O^��F��DyL���W���ٹ���1+��S�E~�湜�z�s�}��S�������j��F\��i�Ӽ�r�bQ�,���i+�*���J�\	��z`���$� �E��ԵQ�Za�!U���8��	j$�`d?���U��H8�Q1Y ��o����V�x�Z8C��_�+��`�qzeu\�{�N���
������n����#U$U�s��[g&�0ǲ�zG�Q3L-帜��i��:x�d��{X�vb��C]�VwY�7����f�!�y.�`�I%�4���l��FSuSn�� �w`�.�h_��ٌ��Q�����2�d������[� u��e�1k�3�c��+}S�O�4�8�e��u�}��']�	k�قB~wN3#,��F�6cE�	�1]��u�D��xί,���D��#wyxd��XD�A��+y[T��p�5%�����E�QS����L�|d�k;m���nI��_W��v�l敉Q�����y
c(�Ea�uD����1OL��V�w�	�s��\m���$���0!��G���D��d�7�)�e(2�:�51�7�=�����o`��*O��l�wm����I(��`A�5F�nX̴.�)f1A��e�_A��#*nW�;��ʹ�@[b�K���@6�Y<����a.K4?��?�%O�h����Hl��;�m����N_Ro�[�QuTMҏu�"��ɰ��6.~�i?Xq�:��.@���+�ߢ�ж:�TI�����9��UH�u��u�$a5,%'��A�s�̊��Q��`���yƧ��^|T�~��L>��(O��ř�}TN�Ǜ�R'�31��\��o��@}Jd��C�K��=���������їq�f0��0=E��
\g0�6�?���5�'�Q�5�5l�o�"��RN�w��l�;=�}B�>a$������{2�uL�7�)�c�5V�X6+�Z��� /�~q9�Ĕ�쪁F���@^�E��f�&O�T��8��Zz�[� @��M'������X�8m�X4��~X�Ï�im�@��^��"�o�46g��%r���NެRO���/&��l�Y�`��l�^/�`������ʚ~�%)�u� -�/t��8 ׼��-/kq0sIW/�-^�.�h����<�����Q.���ϫ��Njg�ue$Hb?���B�F�p qk"Ũc���+~�lR���[Z��^nl"Y�p��
^��cKcs�	8h7�罇�{�v+�MW�\PO����\\��\W�0�cn���+&��ht�J��$ʌt�+�h����~�O,��sd�2B�@-�<b��߻\�15��R��2���r�+t��S[��V�h)�q%�,��V�<p��<��z�����-s��,��B����[ĶQ9]�;�mę��-g��BfT<�}J09ʟ����R��Dx���lk�L҇���t�b���S�yE �%C��'.��� cJ�#���Ƿ��B
W�N�ݥ��V��c�;�_�G�#��y�܅�������C͆���u4�?�{E"DK��fk��W�ҋ'7�E�>5����^{<����!~���T�*L�;�����еؔˍ 4�ĺ%�N������4b�Лe��=��p|N[TQa��f�"s�[>Td֠�x�@17(<|�	�5]>i�;`���UA�C����z ��&!<R���9*h��_|#SV7�7gJB��W*�!M�I��f�)��c��h���|�X��ӅĀ��l�ӷP�/�:Z5������0�6t*���H�F����|�+�"6]��ty��:�좙�qn����lw?X=h��.v�6�� ���v5���j��);�Y��VHs�ʵ��!j�)� G���Qv:j��XwI?�w}B�Z_��Q�������T,PT|���Ƙ�O��S+<z����f�F��
�L�t�b@5a����c��e�c#�&�UYu&y�DZ�#FDKW�#Ȏ���1�956�Û�>-�ٺXH,/6�$�YT=�.���ɛ�7��=|2����???�.�P�u�<!��#q{kF�HWP�c���Pv���gb��|�d*�pX����cZyi�W�=p8ck��K��΍�|	%㧝���>&1���z&m��%�ư\9,Z]�^�&.������7��VĻ���b�`2��kc:�"�2�<�.�E<�V,�%ٺ���!=�㷯�ě�-��:�E�;�,H��@�F��WԼ�����Z�<UL�Ч�f-ǿx��碆��u��G0�^����ĵ��a0c3�#�,��#�e�*rؠ��]���[�e0��p��N���F��$,n>$ʜH4\}��E�j�k��ۓy��N��S�.)��3qU�"�w������En<a��oH�y�V�:mlIkl�k��Q.c�==�=���-��&U�oa:�r�q:��@?�"5�ɠ�U�un�\����N>���]���=�?iO$��,�8��q����A���@ l�6ث>d	% I�I8�a_prr�pXql����u��έ��i�`�ڢ�\��5��`�2s��\�x���C��z����[÷Q^�D{��;�N�8��ip�ʑ��O�!��S?�bV�A�X���IzXג>&/�eK������
���F��6q�ia�k
�W]�2͑}���	�bE��

�bZ�3��^��W��v��%	�x�`�WA�n�q��xdL�&��D}�$r]*dF&�*.J�\�C���T����a��a����@�)�DS<4�=�Q�����s`�-�³����r�%��\ξF-��ᵵߌ}#}��2}'�q���-4��2�&���V���9��n����6����kwM�=O�k��l�Q��'v�$hP�]�wU�x��X.�ZbjW5#ɦt�po����)�3:3B�RSq�nu#�%�]�"i_�r���@�J�9�̎��$�8_Y��V�f�e�þ�5#�(RM(S���פA&y�����
(.�9�d_���K�jp��3�q�� �V���d��g@mdc%�u�#c��b��u�w"^���M��V��F5��6�¤�=Ҙ�,��I{���p�;u�b�Tz��K�L���Uh��ds�O/;ݲ3�e�+�]����BR1o�Jy�.BS�q����������כ�ۚ{$~�횬�~��ڼ�;�Y��Î�hG$��:�*a:�\S�$���&��?s���\^�cQ�6yX�ؿ��O���#�鵷n�)PA�=����CHvo嶞�QZ���"x�]�� ��+z�h�M�[4�?X=�� �dN(m��6�����B5�|�+�ue.f�[�9��C@�j[���Ct��8q������槫~]C�vG�@
��AvO�H����d��3����<*"w��z���]�FW�<���ke���=����%~D�X|�G������E{O���k�N�n9u��`k�����Fٍ߳��_x���&=ڝ�=��,M�9�G�A�8�h;��^z���׏G!�[�7"��6�3xD&<*��⒵U��M�@ީ�$(F��u�m���Y��Vd^ES��s��S� ���3��V<�����ce��Re���Iƅ����?u�_9 c������&w�U�ݺ�}����I��8��vvG�� zo�iUR�w�^2tN,��!��)�u�oO���P�n�P����"D��n)��� ^5�n��3�N�f�,��}�3<yr���b/� �E��g��������sn��D5���E@�dV���4J9�Z��FmG�1!��x�+��H!&qyOq���h;�}�g�ʾ���y�0|�eu��Z���_JE������R59|QxV�&�>�9��fx�ӽ
��,n�G�wq�@X�|����8C�E������L0UsZ[�K�k�R(����j�����!5/ߪ���kA�t�:�Oː��[���:�*�$c)�U}^�$���j]	oZ��h�d���r��Y��&��1Xz�N���l��3RR*����ZO��Y7I�����>TNVO �s��� ���c��[�GT��8x������o�o\=��l��Po�фAB�|zo����g��V��j3���u���<nU�bUd�4~�]��r�W��A�G��,��W�6�2L 'rm���:��)�r���K�g#��&z�*�:=DZws �!5�T5|+U۱@]�Н4�݌��`#l�<js���K`�R�EX�$<�.~/`�}^�y�UƤ>�h�4���c&�e�*�6������ĩc!Y�/P���à)�֣�+;����������
*J�*H,�}���d�ch�₞Z�!/W�K�C�.����V,�ʨ�^ė�� �gi�wv�m�KgY��T��x�:i�����J�����깗mѿf��D>�"��t�0����3���������GP?�c��?�J*tՔm��/�?�d@nz��gC�t&!���<��R��l=���T�"�E��̞X��4H����4 6���=�����"��y�&�hV�W��s��I��x �=���hl�U�Ώi����7���r���yH9q�A*ս��h��G%8o��³��D�#<��~Z�E�Z^pZ�+�G!nh�"�,�t����.�ɏ|C!�H�c\�p�Y)4�ФBCOqq��"��p\#Ѓ���w�����Cis�X�	�����p=�,��}�`��g���f^⩧���--DUBOp��^�"n���zb����澁}���[u��.h���E=Y�c#�Ё�'y�Eq�&�b���xjh����bx� >�)�f���Ѻ,�f�hP�n�:���͋	�S��R�J��1���xۻXݣin1� �TcGc֠0	��H�~�TP�?G�x��0�Y�s��r��Q�},��7���v��_�)�5�
|��x���%R��C>3b�復s���Og�{�R3y�|�b�O �+��>w;yL�(R|Տ.:/~��C���� ��k�BquD�g���}���	���m�jb��4�Qy7��Iۡ*��6�̶Rrj���+{:�s�J�ؔ�d���Q̿P?�}��2 ���H��	\C��y՗ӧ4ڊ��;̓�0�}h�W!���ǧkO9��.�^��i�C����T�Q��ׯY4b`�dT��@��N�\�v؛��:��"�"�8+6��MЫ��4�Pj?��7�v���R߉�~;Jp�'��������Y���E�!D��a��`�<[�d���.4�d)r�k^]��j���QO݂���܄Jz���	��|f����'�ؾ6��_R3ۯ��@qPp�|r�d�}4�?k[�iCgS�&˱���j����"a,@8"��P+���G�3=�g�ݹ�`�_[u[?��+���^�p���1��4���D��c��(4P��X���	�����;
���vI/�t)����n���y15�Ӛ������(�_�{���������]�n�}�r�XA��Q���O`�^j���i�be$�o���	�N��m���r,L�.B��|�8���Ukp���x���O�W��'�mU�@վ%�3wj�=��yV}�n�>�Ʃ��"��W��[u ���X�fi�Kg��u0�w�P���G��SOs��!�lPK�؆���	���~zCZ,��y���HE������d�k'|D��4��u�(r3��?w2�0���������^�o��oi�Q�T�����Ԉ��7Gl[V�4�=Cw�\~�֛z�����t7��o��q=�`ku
wG����0 �)<���?�����F� �������ie<��7�V�q�O,[<jʙ-m����g��v\��Մ��Oa�s:`B����<�6�z���t����ט�9����"I�k�ܺY��N�R.ʡ͔)��Ջ;��;�S��폛;�ۆ��/dW�~���)��
Z�+��0;Nu�kyj�> �0:�K<���>1���)U~�s[�,��ޜ��ϛר��8���x�M��ٯ����8��y#���<�_r#Zw��v(Jp�㯎sM:�ak#W��!O?霔�{�ޖ�:a� �)�	���r`���[[�|���;I��ю��(�'�w��2���0V�/ڛ����P�Cd�%��v������ �G�Y��ϋ����K���,�&�[F��΍B�s���?g�����B���~{���
�g�7��9�F}�a���[ )��V3�F��9��.0��Wɹ��nL,��9�V>bx�y�`�&��?A�v�^������Q��n\4cd��=:�E��SF�>��/�����F�=��un���������Bʄ=d�Xv�㖄�_5��0#w`hyo#а�^H���`����/;���k��P�!��&;�ue�/�C)�� A��K���u�Q�?���,yt$��e�)ʣ�Jk�'���.���_(�b@� ��|T;J�m5�L�����?�uZw9s�o9�������{H�01#uV�����mʤi
[�(`V�%)DF����qҡ��b��"<!��
����`巉r6�Իݔ��:�9�#�
��������W%�+�Ƌ��`6"�d��(�ܩ�d~:���`�
՗�V
h� �XlxVHYEB    a74c    1290]�yjk�^�'G���M��1b��Re�R4���?��!¸G�p��A&��~��fHxL� �X9�K�x�ǉ��齙�VUeEQ���@��1��<��d�=~o���,?W�5�'~ں������l�&nDB5�y�V�?�;���	�|��D��#_�$Wa�@Oq2�~~L���˛�|��8�e�R'@�E�S��H��ox~�PKظ��Y* s�ӿ���=g�1�'�T␿װMN6�dI���%oHŢ%#3y$WV(�Fa��N�Rv��^����Qb?�{�,���5)�_�7Y��)�
S÷��h�Ȋҋ��>�%�z�o���RĮmc�s��d�7���G
�t`�w�׆V�"�Wn� ����+�PI=�K��P�#om�T�99���GN�3�8��58~�h��%X-���&S��]9$w1�Q��1r��=����!N��p�Aw#�G��T)e�o�fn���%��o%^��1��!�X��!�r �i��Sro��������h!ͻ	9���;&��[�N�XcW�l�a�_`|OT�kY����?$�m.������0t���aa�hE��	H�A�f+�����Zh�#�i��~{��~mrQt��%tP3� ������@��(ߣ���Gcr���.j��9�\��")V�D�2{ʓ�j�e���	��}0�x�T8��{l�@?;S3�ڵf�(��%S����z��
�k�E����՜�M
�c��p5�8�2��kC���$�� Ť�;:ጧ��$��Zv++:�^��)�8�n��m��%��n���>{I.���1����s�V�.��hg4�5�5\��_�t���+ދ��:e1Q��������rHi�;����8�*C�"�m�LЕ�\�lu��&���2b�'�wv\���%,���6����������P��a���=e5E�hfL%�_kl�ND�#_�|�ˤk�9�`ì��LC%JB�`Y˺�7�/=�
X����(���{`���5��U$p�'o9��(��oj2C�&�V������yT�_�Ft��,ɗze�?���j��ֲ��B7�=����$���U��
dk�;�D;���rc����ʽ�B�N���nxFe��Z�[��X��6%#�;O�sR5$/�(O;��ŧ٥g'?�˥���~���ְ�s��u��;�R�*��JiM�spK�z��3;����T�����V ,s[Y�����쟶,���Jؔ�j����_��|��W6���ag�r�b����c�8��5Q�<t^ˬ�$�3Ψ0kE��N��"~�,lʷ>@h���V�AYg4�e��f�;`���O,��%���=ë��ؘ��-ޘꀆQ�W[��A\�tF��F���J�	�@8`�4���U!̜R<;Y�&�����w,�O��p+�ER�}�";t��Wn�ń-�nk[���;�=�`%�+/}�ݔ�&ű��Aod*��S����n��|��@| ���-iP�:ݥ�If��õ�	�w�����]�g�2Gsf� ���g@�c]D�M���:rd�k*�ו�uE�d�f*&�5�~��]|	;>Y܍�%/Z��P���KK�i툎:���/�o�|M 8�+��a��r��ߴVC����MCH�n��)����c��-{T{.�}����%�Ie����+	\��)���tqEB�e��r&��2Q-`����k	{
։'�%��ۮI]`����x]}�a����H��#��է@�v��U��\AN��M�G�ʎu�$Z����r���wXS\��R�[���-��T[�M9>��kc�*`���<���X|X��B��n�V'd�<���@�2��(��:�e^�����Y�ޣy�ϧ�=��N4�|c�̓��aV��"���U91��D�7�����ٿ[�$�זN@>��h4ڪ�|��W�~�Q5�g!��y2���嫅�����[>�2��+a�|��p$�p/헚`���D���6��9�3)�'�c@0���GF�1v�\}Z��p�!N;�M)��3��2����8�P s�l���>t>M�+Q�~�NC_8r�S	z4��'�C;]4E��ј�r�����%z}�#�̎�f*vRMq��&� �,��N�)�'9���h�<Ё��Fj�
yn���R,61#�zI�����,=msf�m}]nv#�&�N��4����`��R�}��E�a�;�� �����y�P��h�Cu{"�`3z�����ڢ��ݥ���/n�����/�4�kj/��Dӷ|i� ��������%Z}ނ�G�ܪ|��S��6�W����P��6*���d��,�-��J
 Z���j�
-���z0�%�n�/� ���G��"�.�l)Bu�ݻX[*rYG��]^�8�"Z("�!�g[��;�t��ľ2JkC���~�vX�ë���j�X/�E���}p�z�n��9��w.O�l!d|�L_���X�<�7DFE+�S�Ǽ�U�[b�i�F��^ʊ��["D�I���~㒽������g����Y��>ғ�q�B�����QJ�\z��M�"�G�N���f�S[o@�%W�~�	��_�E��fd��_�M>�+���Y�o�J��B��y8�V%3��)�u�c��@�~�_��O�Ώ��bOP��nU\����x��>�&فyaMH�{�-z&��\�}J�Qf=�� �� +��O6�f�j��O3j��xZ�b�&1��9��������j��~81$_���o��G�k�<�q��C�RP]�̽����X�L�O�W��P�"�������Iʶ�Tqk���}��u��N� ��&ƤM&�5kP���B(gZ��"*x'�W�QҘs�Io&�mL��}�^&`��������U���Ac�b��:�͙X�P��*�A�T�JY�8�3�Y�,�]����Ş�o�	�6� E���i�6�8�����[�t"�����g�SO�z>�~�׾[�G
�v\�6�1��y�rW��ڊ�!�(���#&��V�>fI	�w�- �3�̹��L$tt���ii�r��D�_��5�C�w�{%1�W9	_�$YhF�X��2$e���ax��1�G�"h!��}��1��
�$HN:��
uX�y���}9�g4n6���9�*`㝊��7ʯP���8�fԌ�P��|�ĝ	�acp\a�"�?�q�u��
 &vH�&d��.%�3�O(~�Y`����{���cd��>#(�ůb5|��b���bd�D5ãC�I,l�ӕ�@=�1\2<�2nܑL��"��y���M�2^0k�t�!��5ƎV� ��l�m���F�Ǹ�zCu������tH�)y$�e�=Wl[�[UC�yiASXi
u��\���{*0Ro8��q��'B��A�I���1en�qH��%������SvmrJ}��I��7�F�$ﺹ_�kW[�~��z�./.d�E'�'��NpN���+4^d�W�J��b0N}r������(rA�
�hy.���
���!�j����8	X~'c�#�<l��G���׫n�v��n�c�6X�y�s�l:�G֨���ƭ[��A��#!�]yų@���$��LȽ_X�-�����|~դ�*��ޫx�5�t�A�Usl譆�=^�{�#9�"��c����H���.�]��,	�J<��8�i\��q��L��=R��͗ѽ�B&}m�Gێ,NJ��Um�vܖ�>���_�cI.G^/�$�X�t~ ��z�YG�o���F��å�8>��Y�����^�O�	Q�kj�Xs˘eZ�� ���:^�.��&��Zw���M������b���}l��u�~^>�o
q˖����=sH���S
pöI�(+�Pڙھ��寭�v�Kt6�D���Pj;O��_j@'�/0<��ʛ[�4��H� �;��Zf�^7�T��4)|�y-eu�N;�l`E�0�#\Q�_7��UrJYq�|��K�Ȩ�݉�xp�����d�����������L�[�(Q��.P�] �b"������w/�z��sU�[�m�3(u�[�j�w�b����p񆪈 ǽ�����t֭����?sr�yh��G�j]�ںn0�s��_��&c�]�_�s!�n�m���r��f=ǜ�S�q����W�S:A@Bec'�V"��9��>�����Z/+1{�l\'��n�s!%��4B,m̨�Q��lr�x:�௻I��wf#W՝'�oQ`�%؂�����v���7%X����� a=w��^�x����ֿ������Y��f!�y�5�)��	>ɨ�cUv>�$ɛ��~Fas����y[����;�r��ݟ��s��}ڔ0mȝ�&�`�Q�����q��_;�@��/0~��KȌ�f&��E> VWng^ZF�$�(�Cf|e"J$j�X�G��2�é?���H`�[������|tt~S\�k��py(05K�j�����M��3��nZ���m�����M��N��L�����*���K�za۫�dМ������'T���j�H�}�eE��!QX�{O�*�$�e>��bf�״�\����̻7�<���r��硲ލ�]�*B}�ҙ��UF��B����38�d!�Q��<��G�+%���.³�-�3y3����@WŚ��`g2�Ah>��>wIaz��=GW�