XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^�{���p,N˘��CETG���U�d
��і��dD��C����[}���n�N7�W+�^�3���F�B:�����AנK�~�����36"~�,$.�]��C�	���$r�	za�u5V�x@MK�AI�2Y*�i������W�뜃+�a
���!>d��9����)��69��q^�!��C�B����G������d�](aFV{l�<|-=��M���D����?k��c�S�A;T��sLB����hKD���Yˆu�1���N��$`a+<��٥Ϝ:=3~h���v�m���L�Uj��	�~al�?��cP$Uu����Q�y)����nR���ҡB�x�*�ƅ$i=5+|����%�������*�F�Q�̆sB��[>��"2F_����x^�! Qˤ27�㰎��o!*����w̲��󭫡+::{}k�z�B�`g���� ���+�p�5 ��yV�{��)��>�t��RymF��?�м@���&�`ʄ�^=f���m��`8z�6o���A�C���0��tK|��!��O�鞯�M#�8*Q~�h�Y�^�.�4�6�y?�آÒ����";�?Ķ����J������#0/��rO��_���P��)��_��9�����p�t�3&���5�%�B�������M�X�v�C�[�L�~����س-�(#t��V�������:��[��Jg)LV?�a����bZ�j!C�=ۆ�5a�pV�N��XlxVHYEB    302e     c70�q{�"0��h�ڧ��������Y�ڄGۥy6 �{�n�Ս�����< Y�V_����ɢ����9���(TGl�u_~�����6v������0�3m���mʳ��]�e|��%̟���	DC��*���s$c&�^�Q�d^���Hyg`�Vr�"GuF�_�e!���t_�^8�D6��qtg�����Z�(*z�h���s��n��5x�Z�/Ct��r�9�~�Gi%���?;eR�����]�������h���f>��K����ad� 8Z��5B<��.��B��F�e؅�hX��gy�e�����f�]T{�d���IRɆ�ǧYt�
<�ʈ�45g�������{��!����WKv��_j��K�ުɢ�e������L�^�I���fd�C�-n-o`��(e9(�_�a���(VU�38#��˜g�ߛM���� �f�o4r6�� �9�$�boIq�YX���AJ>����:��aĊ��#���؋���\��N(���"r�Su����+���{� �7�in�����P�7�q�����V"���k�箿v�~��-C��vB���+�e(�	b$9��� o���T������4닽�״����-����������cݷdnζ�;a���������Kw��/���M&���	�t�w�o9?Vl���Xٛ���k]����ޮ*w(|aH�!��9�%gKB�=�|^��Э�0�$y֋�Lfus�c,��-y�_޺�Z�u.��.3��1��u�k��ٝ��K�w��C�7��Q��7�����.�-�3�-D�Z�b��Ǟ38O��8�����/�V��8��Wn�ד���Z⸱Un`���X��,�K�۵R+[����9� ����=��2�M��	)��+:�&�O�	��+�\�D9I��G1�,��v��n8K�[�Ԃ�I7~o�(Ő���S��>�/;"�a�g�f��p*�u�6$g�=�ݢv!�J�C���M%t�of�?��9���!�u-	����#T�^~�
 �6��h�����c����q�R�0�`��b��4�J��W�e�9 e�gfa�='hY.�s�������:��);LU" .�?.�]%Ha_�D�q�I��:�s�M�J��o������h�ZM����	p�Ճ�D3����ɤ�X}_���p���T�]��G~�<g.A�	�7����B���g���>��?M��3��ЃQ��=!50:[�2	G4K�n0��i��F���� x�[iZ�}~5�.|�K�#D�ޚ\�ᖃcd��H~�!��\O4|�ƕFJX�T�Qp)BI�7��8@�G# �z����f���bv���F��Q����X�2�ތ��J��l�s"��g�K<��Bj̼����g�(Qo����_�l$��-a6̙�X4��P�Z��N>$�J���%P��ʟ�*@�ڜ�Ӕ{H*�Z�&��q���<��v����S�u�)�R�'�n�5�K��}��6;N��cS��������d\�	���A��Ve�g��� ��C
�yr�Y+�X� ��sM���&v��TM���=^�d8Z]��bT$�"�2$�q�T�{:�*�أ�H
m���:��x��(���@�Kf�8~�/�5�i�f����� ���ٟ8ˌ]�g\��
Cba0� ��8(�$���s՗>7m�
]�������+��0 {�\�X�l�]�X��}�*b	�KH��R\�A.^���s�+w�y�׬4u6����&�8'O��B�1��6s�c�$�� �����ߨ�2�OX�p�A�X<�����%����yF&���Q@�o��j�*�*��U���b�:!`z@��1�I�/����t�?�����W�\��3�E�Ei����*�3I�b�q�%6���0��+��F- a4����#y�=��HN�F��˗�cp_�0 �L.k4�f�����O$�Ј��u�m�h���"��C�=]�2�����D��c�8=����]��q(29"S�9ia�7Cu9��p�����@�1n+�t&:zB�7�0b�ł��|2�:!�Z[�j���1<�I )�F
�{�2!���2,�Dǘ�՘4��<<�=]����UV��'��󽩚B��2��Zr�`'�WD�7�C$�Y����6�\����R�h�؎�۬S=k��#W��g��A�ɥ�ЁB/��m���6�n'�	I�+ߌ	�Kl���V�+�a�LDP����� �|�(�6�ϛ��$Nĸ�Z[h�02�_74gjO�]�m-t�2n�l�z�*�u���l�VQ��D�!|�h豼{�J$����(��75�n_ Yw�+9�U�E}԰�|�A!��%�"���o٧�<H�H�4��&�q!2���F�5IuÆ�40jH��nfM�D1�`s��7�����]��|��rO�}9K<�p�0�B���+jW��L��l6@/�#~���gUѺ��M���f���	�Y�"�(�j3�Jw�2dEC�bKܡ�Ba��ru��囌�8�,��޾���:��*�tC߯�#32Ts�а)EA��v�àż�֤�C�e~ʦ�Yf�^e
.脜,�J)*\�X��4ĭY�����i��USZ��s�U#�#�,NX_0���_��-���3����P�tl�8N����DE�=X�%�����~���0����F�L�}Kd>_�d�����`�twfЫs������%+C=gǜX��8uO�����,�8��X��B�u�8�B��Ud�� =/�/q3UwQ��E�,k_�!T�/N)g)�B���X5y@ে��K��"�9��1��.�A��/���j�R��@{������m��g��8�z�m}0m�����J���2��!U����	�����+$^˿�Id2_��]��셫�yNǛ��e�m�R3��d��7l�Q�ǉ��/�17G����S�~x;>y���U����Y�0t�vqɧ5N>\A���v~\�=(&�v����ȹJR8]�)�WS'A����<U~��f�%6������Jh�H S�ٝ�rӋ0����&b�C���=fJɛ�!s���b�W������F�.�fA��t\���e�A>�{��ԧx����87i