XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y�;��!���Xz�7��s��ͨ�+�s<K>�o7�9m����!�[��~X7�X���K�/e�a_�����5�S
F������=�8�
sN�lH^'B|����z�ɹx��0t ��B��ݒ�H;O��g�B��������cH���ei�{rf��;1hxrb}��PaF�S.��p���X���.�;�}�fd��z��δ���a�V�iL'�f��)�|�VN �����)�c�\��c=h��t��f����Aؔ�Hj���[nc��<�W�XT;Gh�ڞ��n�R� 2y٫�T�����)љ4���p��ڃ�MB�UX�;�?�%���35)�p8ɩ��c2T���3�F)���KOi��0�:{���Ԣ	�l�xkz��`3-^��v��L��n�n����l��/����?�c�g=�����,�Xd�a��ר2Q;i�Jʒ���St���DY$u-�>�����pZ�&�����I��R��2����m���i�"NV���e�&~��\_1*��i.��E$��>�wƁ�7��>�p�`�4���>|Ѳϊ_�MS8C4�!	s(�n_��G渨A���B��U�1��$�3M�Fwo��OWxZ��#C�/��6	����c;z"Ak��¥�&A��J�>f�(�\x��
��5�dz��ﲖf$~�����1�f�p4H��\�~�T�,��'d{O�i����%�^4�2ESASa���v+qʫp_���	�N�$�նXlxVHYEB    160d     7d0�"d�;�R\xv4�~��n����R��DQ��O�ؙF��r��Ti�%B�����+�L��8F(��|AF"��l��*bL�kS���H�t��5dc��o!��$� gv���v��7^f���lTS���3lgXܾ��6���U��^ZR`}�Zy��u�&@�t+�Zn Ձ�C�/]坈�(%e&�K4�݃��oR+r4���?����qn��J���7h�D��_���eC1�֍<٨�/r!�æ��ǋM��T��Dׄ8�C�2�FM��!�OG8����i���yg�5��d���5�z�H�(җc�:n�zm�nQտ?Q$�iU�"����h��AK��#T���Gz�+���@�jx[���K$5����ϒi���IM.'�q�^�ץ��R���TV&G�۟�9N��G�����\;�)�5c@?�I�K|6�Iy$5��3Ю�����}U��B�@���T��t)NO��9�:��x�S�]ܞ�n+�3����)���	Qkʘ��Z�����|ʷN���A3�&�a�����-H��m��ߕ���%������$��_�m8�$��w{6�	�6��ԇf�� ��G���H:�AVA���5x��v�r����kY���S��>�w,���2���,t����A��~�Js�����|�o���2�3;8kF-q�i�Ԣ��1u��>��d�y���T�Q`��\�#ɟ��`�!��N*�AN���<I���95	a�8D��X��py�zGlIM�=��c�ս%7�Y���.-��fQ���	׃�=�,�Wu��Ą#�(�P_��]F։�d�;�+՞2QD��x���E�P�ˌ<�<cs�J��>C�ҕ��-����a��?9�� �_8�Yvc9�:^�_�XA��3~�Z�77G�"C�8�����vV�)*zK����%Y�3%0=�v	��
9�����g���t&�fl��ۭ�ׯ��Q�c����Z���֋'VH!^�� .ɸ��@,��O��@�Ǩb9�eV��[@ʬF�3��;6[d�S�ǘ#��?5�&_�����`s恲k�H�U�P�a���3!��-S��<ݜ���w�W����+������s@�Q-FKcF�{�R�7ˊ]�䷠��YN�Zk�4J*C����3�Y9�>�{8͖���N���G�9y�Z��(��.�[�i�,����d�ʷ��f��dSp���g�Qu��(�3	�wԄ�R�O��4�MN��4���#aS�'�B�έ�#[�0eS3H:��LƏCQHP��>��y���9+0�ۧysA��3� \T28_x�������������j@%�*�p��>Ъ3hi���E�M�5j�����:![�d��rӱ2%E����x���h^G��e�1y,���T�6s��(�k/���?'�g�Ԯ�_��e��H<�tإe��͂�."�i��˥�C�����#ѐ߬��X�"�2?��I^�oyU������i=�T���N�{��'�ju>�^ugY���ư+��χqB�og(���Ϝ��<�6#�_Z:s�����zN��bFYL�s0K? �]d?*09MJ7]������{�v��V�[@Wѻ�s)�~���.AWF�c����9ԝ\�9��r��L�9�|�C^yD^J��s_��J���^�/pu�VĘ�_�z8ϖ�Z����0�V�;]
�G��=t+�9G ��A!�?�v�Xl�mkt��H�z[_�֔Y����(�(	��]9�i��V���o+�F�C�x�ϕw�x����_H�s�53yU%�\��e�*ŉ��o��U_�J�7j�.��.�"ڨ����)[k�c��G~��,�~���V�cA�tl�) �n)��Z���k�^�����l�01d�L�=�Ps�1�(zk�q��n�@̝�l�%5��E���[" �:���oڹU��~�_�&�,�ڌ޸���Wke22yb[q�YH��_�