XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Sdc�C���|4�K+W7`-ƲP.�j{�}�p��Ә��c� |��e�W���ř�B��:�������Mw�j/�'^��;9La&�")@):-��t�KO6���"�lC"�S���4�XC��b�r���L�4����?�+m�~_!��$�^�J�[C:1��z��a�һSr�??�e��(8Ix�D��v��)��m{�%Wt��+�9=�8�e �������)aD}\��P�ג�k�����g�Q`�5�M}�!�>�of��/W䫮T�~�S�xM�bu�J.�*{�2\?}�be��
fn�f�u���L�a�I��q��x����h���ލ+��:N0��c<�bö�/��;�{��D�|��cJ�'�	ۗE6ZH�7�n��Ҏ���mQ���HL�M��H�:͕1���(�tcN�����k��O����M�]��}����/̛}��l|�UV|�I�~pշл�����dN+��d���w�tԗ�$EP��Me��*巆�W #
����`{v�JI�`�_[ ���Q�Jn���@���h��+�ĥ�V�v&� ƍ{[>���B�5��X\"�R*�t�fI8���人2�,�HB٣E�G�&{�KX8O�I���]���0G 9ڪ�ۧ��Gw���ũ��l\�褡fw�KlV_k��ƞ��� ��q�`[�����p��.8��}���{	Z����@���癯R��A�b̰��jF���rXlxVHYEB    4089     e40{=/U���AU����ou�Q�g	d��]�q"\(���#�j��!����p+��<òɵ�H��|R���m���\�G���dN�х 1��;���V`h��Y������㪷
�� ��� �1��͔�n��G�K�G�h���
�	�2���K�}����TDu��d?K)xu���/�^��S�C�;���kN���P��>3p;S����33"���?��e6[!��Ϊz/-Q��`-�9e$dH�&�B[��-��4`3�sʤkh��8n+�� 9p勧t��	��Z�햾SιT>p7=������g����Cj�U��?B���e�O��8�W��=v�=��� �C��7cqp��8s[v"´v�����m�����l��"�O%N_e�P���C�t!�py��N��/��^���ּ/V��M��-��:��Ѡ���Lk���q��g'�p�ٽ��j�'y�H���9�lTG9l�4ۯ^���eR���C���TL��w��f�����= \!�<�M(nw�Q?�:cLU�1H��I���}�)f�ͯ>Dp;aKFIxh�z�1�B�1�lFpaf�`�{���.����u�!(.t	PU�G>:Ӭ}Q�Y��6����!��3��c�`�CqE͈���B(���1���ڨL��ht�����\��~�|T
f�nK�+��+�88�J�PWղ6ĝD�\�Z��	h��Ow��o78��O'[�R*Ȭb�X�� ~�.�<��ĩ���n�����>%=zy?��Wb�܍���.���|^���>cm��a�#� Y�Y���XM������5��A��G�hO�Q���2���y<J�TN���+�ߺ��XxQ��j7��N�n���u>2S*g=}6L�L�)ۊxt��i;!J83�ƭ(n��Y��P�g��-:;.Js�6~F���\Nްz����b)م�I���$���\P{a�M�l�1�!/��!^:N�G&CÓX]��+�7��r��جٲ���1�k�h�%�*o��xo<���k���gG��A���`��k"�7�t��Qt��	�gY��=�4�DC��kzwӧgᄊ�ka��Q����!Ø�@HK���T�� `�W^Z����3!Z�����tH���d:fp|i��li�j�2����ED�����8�S죂2�9�[�ꟹӐ9&��A�"nʒ��{��N����l+	[�i#^TL��̊�+�!��]e��m3F����[���ƪ�:�	�T�U�?�|��C���-GB�͝�������ouc' �n��(�A�}���_N�_3A���{�U7dg�e/����/'���r��d�1@Qd#�R�����ߩ�d�-��F��V��o�m�m+y���[��Y�-s��QV�>�U��P�6?~G(T_v��!1�L��_W�T���~��4�A�;0(`ϭ ^�8��N�Sa�LZ7�qsq5�j�Z���ogX?�Fs�t�j��
E�+��2]4�"۱�날�����b�G��p4�co}T��J�4�������$�C��_)���rw�*���~
���?�<İ�c�|�=���
.�Ϣ��O�`��Ϊ���H�����(�0�4<�s�r��g�:��1�����I�	Vo����2rߞr�����G�y����@f��p~�ם7CF��>:�L8;{9$�W&�/\�؜xA{��sA{8�� ��[��>��=+s�>QP�`)��!����e?+��:�''u�=㷠{|c;@�}F��m��(Aʤ�N��ގU�*{f��+W���&��,�6�­b����5��\oZ�S2����{��Zk� �6Km6�dm�	1�T���5s7r�-�}�z9����G��i�'3�;o���8��\��
����|C5���p��#=���ώ;�&�CZA��	�V�W場�M߼{���C�x�.j��4w�ķ0^lJ��]7�PҼ�}��˚�`�9XUOᶢ�`q)��mж�e����8�mC�G�gdu��ғ`���wv�(��汣,�=s����ig��Ex�����h�3۲�V��P%�Y ��  �2<�����u�@��[$�Y�.)���Yj@��:�p�x�g�������\��ُx`�Ry�̍����9�ƣ_׷k�楘��O�m8�%�	&ch0N����q��zR�	��+��F'�I�����Hx��?(t�b}����HK��C��R �$��9�J�:�ꆦ��2�Z`����Ѩ�B�6)����N�_b�8@����_�pZ����f��'�c�.���.EQ>L_��FA�j2��v�W{���v�qSGC������(����R��d�����E%�/����(U����U���Q5~��Vr���>J��.-aBL�h�W�H���]MC�EE��7:S�;`-:(�t�9^�)����!F��>%Qc�Zخ�l?>�q��	yQv������pNV�f�$P�16�yU�������qo�����/+J;������^��;���<oh$+�� ���:��i��6��#�=���~����u���� �f�]�D��R͖Ռ��.l�I�@dv�SS�KZ�4�Z�r���f�\�&�<��:�����;�}0�%'�%W�6�hٸ�"�b��Iv�'i�m!K�B� F1f ��f(M�oF̼m�E90��.UV3�ӥ�# J䚉(	�E��RL �/�X�6��}B��I��U��Fw���h0��c�Δ�~����&�%�jzT�.ُ���Uy5-M��:��(�2�;Zi{*�ZJ	߱�`�g�����t\���H"X\w\	�־�j4.���9pѲ��(*�Jw��{�a�C!F7�~�ۉVP��T�2SL}#V��uC�!���M�:o�8,�4�_k+z�@�t�*�q��80+�N8�nX��7���<X3�p�<�n��.���-<+m�d5�~��DGe��ɹ��_�x�0���it/@"���W<F�"T��ؾ���iPM����r�	�!lD��O�7��0�m�f�f��dc��b��/���ً�<N.XL�n��C����&��<� 
�uq<��B����ЎW���ts��"���`r�.�j����G��(*4�w����j�6�n쯵zg�-�ˇ�X����5TGY[%��.Of���ë���P�F�Ь�K���:�	�*wu^��ͭuU�!,As30"�><1��X�s�#a}���Eժ�n5i�ɍ��rt��u��ƽ���=��������A���j!z�Z�AC�ֽI�pΰ(��n���b�i�0Z����a2�5�xV@oB�0��,c�_W,i����o�Ma�sb��2 ���祪��G���-zx�
�E��"�_�"4|��X��}>?��v��b�j5x�iFl��K\�t�������r_��u���hu_���d�\ec1�b9��,g�w�.����'-O��� e�`�S��BGC�!Kb����OI�̾'N�y*%n��
2�n�7'� p'��`gp	�S�"�?/��$�7l���p$�R���WqJ*�T�!��+�] �`; ��7��ڭ'!�"��B��