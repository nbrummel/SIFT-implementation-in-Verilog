XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��qCz��{�.&�%��~4{; 6�_��?�e�:��p����P����9��I�f��\z��{Qr�^҈'Vb����Q��|�����vF<�V"�P�ڙ�i�=��O��'J)�a��!Gj�|aʪ�)X�o�9 E#`�E]�w�\B��=�1��+��D�ugݤ�f��z��gM�2��g������j��'����Ut���~E�2��*'"_�1��o�x�xa��";�*�k�?Q���`%���(��G:�w_�=�<'��H�v��ϖ۰m��m���L(CNh�"�n��E�����is,�Y�/t�!���%�����bdYk���������݅��1��Qk�%
'O4�E\��2�n�l?�7Z�!��1N�����.�o��W+n��o�\:s�we����rs��q����Ydt��w� V�/D/��x��5��>|Σ��}�^I�@
��g;p�,�秕}��-����KUv�/����%�4�e��5J�T˂L���G�4Ҧ�k�=wr���$K���嬛���@�^)i���{�<X���nn��O�t4g��o�_`%z��d��������;����`˲in��܋N��Y�]|)��^���:-}���{I�˿d����U�XKzߝ��Q����wD��9}�$��)�8e�6)a�ɿa`hX<TY�Ǐ,��]�T��T���h[d=~�iHD���`��60U�o��//��� �g_�m���!o1����fP�o8XlxVHYEB    1ce4     9e0�@W�����2Bce#{���8�	;qx���r���.����z�9cēG#/Ε���;��\Ə��bb��(lu��G 4�ʚrl$��w.�Ae�n}�^9F� 2�.��R��q���zkϳ��.y's7�ɇzGϕ���<�mfY�E�[=�{�c�o��J�]��a|�g HDF9��uPD� 7�d5����!�<`��9�;���+|�U"ڟ��S�e��T�$D3�E_M/[�<uݼ	iA�Ha^J�P��R�ȝs���/k䏇:��D&��l�)lC;���/ڌn�IC~�w�w"���At���0�̌��Oo���!��N��9*K��u��gcNE� $"g4^����I�ҷk�ن��9[��O����7�+pVP,vF��h�_�关(��V�	��?�%�~��� t��߆������6�׵bqUߴ$�y�4�W�E�-��@��<��P,6[h+�BءRycK�7�R#6��n1*z,+%h�i.���n��BH�$�&� �#zR�r�]U���n_DU�pڔfU*��w�ц��az(�l� �0
$�������c�+2H�h	zp�j5�7βG&(��P��uND��� �h���{4}�3��\�^� fU�7VN u��>{�tf��/���m2���n��)��le&�� '�È��� :��ŚD�w>u���$xP�n�G"��C�7�y�xFAH6�ᇽ���yL/������<�[B#��,�X���m�r���/ߔcH��4��c���=�H:�A����7g��WbG�N�h�O����΁k2�"N�Fv�EK���N4v��Hh���(u��^ <����st7$�
�m���	�3�y��L�G,7�qrٔ�:_�C! �H(�%�]���Y��u$�_K\FT�r�ŷ��yBV���.�/������O�v٦R�胆k:�7@ur�b�bh���el?��e���{Am3�^Mx�A���:��% >�`��׆��iF��/��k��J��אH2���uJ��c�נڵ^��p�A��I	Miլ';���fX�=����~�O)�0���N�J�^�9��(���G�M���|5u|(O��\���n؞Yxm�O��1=������n�;�d�n��60�0��v���l���c�`����H�ffK#hb��s������D<�!�[&��0��jR��)���Y{1�RL
A5!�?�w��/��6�{�m�d�lv���,����N���~�Qj4��Q��C���C�7H��m�C`1f��Ǥۤ):��b��Q�F�3Chճ��Ы
%�0P6��FW��<2w7���G���M׽N��#?Z�Mo2��H/x���_{#<g�1����l��~Ÿݲ1A?��hD��W��ߔ�_�I��f:��#�@���C!NP�nE��H�~$�{*#�2UW�h�秞o�Aã��`��!�k��&�qF�)d��9��4'�d~t.�(����&�>9�w6rX�ח٧�Rw�!y�S��
2�H�-QY��'(���< �m��Z|Ʋ��*����ȧ�@?�Ǝ�z�Q]#���y�-Ħ=��iY�GH����O�yZ�mD2I���[�]����n�8!浸�B)4h34(��!
��Ôϣ�i0�1{Ex;��^k�n~`X.*U��b�͐�������E��UuT�u�D`�Àg�{4FBm���I2%���FJ����"^�2S������7��0�=���\z�d:�|	�|����<�TW~5A��,�,�%T�T7J��r��z��Б˥��n���n��;�����9�\�Uu����Cf���g�|o��Ds��g��[B�uG9'o�������4ݼꎺs)�@��	M�L��!]z�q/%��C�S��B��k�E1-��'-t��+��J���J�N�L�M��
���x��z�r4��� ���Jv%�U6ϙ�8��K.��k.���8ױ��ԴP�k_)��~����l��@3w����e��DӜ5�f<�g���(�V<[������kǧf+w���DF͙f��CAv�Ei='�Q��wȳs�iҢ�����d����ń�+Sa�yFh���
X�k�r2P+'� ̬.G<�5�G&��Ч?N'�)w��!Z�5�箫���daB�����%tp| w�����شC��c%Uӱ
�"6��*W)Ci㹏�	y\���y0���Ea� �.>З8��F�#n�_��y5ր��������Cw����.�!��z"�j4�F�6~1�4��Q��P�}X��v��U|���yh@p�ÂI��z}�8'�';�)�S$	X���W��ER��)��}4t��[*E$�� K��tg��qί�_��$Q5��$s6�Uh���Q�r�|9�Q��GT�G�l��۫_$6&�I��
q��+o�t�O�J�f�<YL'�^j=���=6���p�x�8���e
�H���w;�����0���U�|��r