XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��iHK"_���$��wG�W��F+)bc�_k`-��8q����);�j����&����ٗ�,�����A�B�yJR �'�A�_>X����k,	M�:��M���Ն��F+a�[�Z��X"�{�IeT$�}v# ��{��?��X�U�u�x/$xr�<�˛��b���aT���T�=0�/���ЫDidX�X+��5�k9�Tѿ�����f5�ɂ�)�YwNVg-.΢�L�Ӏx�/�zډ
��{����h��8�8��x.͡~f��"ˡ�_r�C6��3��#�u���z�׻���yy):
��6�	��R:��5�Swe{W��;��b;�d��ًa�@ƗC�f�H����6�ؚ.��ۀ�ȇNy����ن{l��3	4|��V<�=W�Ux������*[δj��Lg���#)T����J���t�,^3,ƞ�g#���o�iVI(��[Ǖ���J�ch��yW딞����M��l��mR��+f�o��k�`�Z�Im���G����IY��4�t<U2�����I`����IB��P��Т^�Xc�w�B�K_��1�Y�ǜ��\� ;��;oay�_�� G�F�}q��G߷��u���';�lǛ&�(�[>c�|*uX�c�u?v���=�`])G���\*i���
#��h���Z*��&f��g�C8Y��z����-�MV˅�whFs���>)\�n�bw��d��|S����۽�%�3XlxVHYEB    77d6    16f0OsE8p<��z;U��=~"էo���a+s�a��4�zk�vQK�2�k��pè ��2IukP���QO�,���I	���_jj��\J� ��jSv��p��������4=߸t�Հ?0���)�Zϊ(N�&��8�,	����BVf`��]gur�T"_<7�!�`�F���o�� פj9F_d�ڃ���wv���6i���;��<ϋ�E�\7��S���-#�,w����D�b�U���i H:� _¥�F�P9���m���I�3OQ��@jQ��u1�.]v#7
��a�M�&R�!(�?�ͱX=�u_�Ǒ��{�HV���1Oe�Å�����w�q��p�G��!R��͂LQ�q��s"R)r̳V65�.���(�!��־g?u�@�(~��;M��M XJ�n6"��HD��ƋՂ=&�K�R��tjL���OH�X�J�<mT����Ne&��Mv/�����zc��I�-s�AF�M�	�e~2��q[ ��c�8ȹ����d�,���^�Di����d��4������GH+tQ���Ԫ_G$dW�f���� >���~�SH��(���j�W�+�d�ęL��k�[�g>�f��|ڋV�k��P����E�4�
��G}����ιƇ��m��}�|���`��X��{C������d��hY
����.��Q�&v��@k�נ$����o�jn:�8�8��1���T��v��g���O��Vu��g��9�{�V}�Wx�(	�R��̅ �gJ  = ����F�F8tP<1��.��gP�gm8�7�ͽëf�7�� �*�aP�_
�>�g����1��;��Zm؛G��#�3��7��z�D﷨uEF]��v1��IU�;���<2TR�ٗ"�s�Ȍ�M`޲��}��i$��Ts�(ԟp�+
6��M^�i��<��#��*��G	�������$�=���[@�RPs�Nǵ�1�i14��:2���A��J�Y�%q^���R�l�8*_
����p��:X��A���� �Iz�3"�<���'�.ȭB
B��л���l�J%�F0 ���a��>w#eE'�R�T$�M�∝���i����p�m�ɇ֘�n�I*����_�a�\1�%�PG�њ<�1%���OQ&��;���h���܊|���;p $����鄏Ĭ����e��f�yl�ǯs����^�4Q��v[Չ��£�Ⱦ���+u�j��#A�j	;O�A����22�'���!o�ܓ��[ ����n�M��$����ώPϼD!rsT|��i�v�*�V-�{�)+� ���ؑ&52�U���O� M?��o� ��]����fb��T�^L�f�(M����k�fuq�V�t
 y���1�s�2&��:�F�V��ό.7���u�s�@��E��M�����Og�θ�4{�k-�dk϶m��[~Wq�4ofO6:�� &*�d�SB䚝n��r��y�K���Q�5ȼ����#����v������8 'F%eP�V�y�n+7ǭ��b��Y�goAS�6o���ffâ�(+��޻�04��j�(l�;*�݂��7��]tY�Jܴ�q�^ P�ؙ��Q �Z���,(�(O���&���SI�x����ܛ���}s}%�]��W�eB��2b��I��z.B���}]Y��}��}�k���Y������y�\�}��1P��H4�_�}����U�QڅM?	�X�f��([u��T�19[R��cK��<��Е36
J:��1Kٻ-�W`����@���'�z���t�1-�Z�:�&����d�q����~L�����S���nɃ�����wD�w%^�����"gQ���%$���P���A�
�2�gB�T�2N�PݿI�G'ȳT��g���gDbb!Ofp3߭ĉ�]�4C�h<-��v}I|�'!�Iu#���1�s��:ː�v���.�ބ���w����i�\!���VCC.��W�ß3�g���5�MN��M���L����	-vŽ��@���D^�[`娫9�z��m���w�y�\�n�0f9R@�C��[���sw:;%�U^*���⅝���b��Nk�B�F��G�����!��$�Ds�,�Q�6>��zbX���	,\���_��Mv˲��Rρ5�a|a����A�O����GU��[�#r�_{�ВN�|�����΄|�k��;�w�.�$K� ����AC�TiL�Yj@��4��he�f�����K=Nn`��+ˬjI:��~g�E�E)(�n���C��z>є�D:`[��l�������Y�p ��îV����|���:��sd.��7G�556�������Am�Q^�J�tN�$�2���Ƥ�"Cmc�Edct��F�����K�8���>��ǧ�M�m�$�4'����]v�w~i\���ߓV�nm<M����������\��>Ǻ�k��������"4��xnK�C�ںHc����R��	³�]ƒ�qr�a���)9�2f��Z��b"�����Q%z��	����r�#5H�"�u�)�t�-o����*%Q�U��m�Hz�KF�e�F�g��[y`�T�y�_����NG�h�~�I^o�������>��ʡFc,Io�4	�5��yM�H����<4��� �h=3N��6w�?���޾���&[?M�vG��9�s\W��X����v�ZhWj8% D>�_���o�����5������\uq%�!b�L���j0�%&�~�G\��B�	'5p����DUB��4D#� :�c��{z���`/�|��c���
�Q���rFTg� ���^|�[Ʈ�n(�����y�a�m��m0��������2����۶6<&߳C�|��PF�Y�5R��B�l�W��+���$��a��G����_�}4���0\�!����v}�g
B3>kKhƦ��a�R>PJ���Ύ�q���6����N��v)� (����uE��^t�9an�,涡"ay���&��%�4�z�/%
W=U�����ƺ�9-���S�~3�K�����*j�#������c��<��`�<- ~�UO���2��7�T��qJ��3�<�Y٬��݀\-���Bi۷Ü8ez��d�o�Q�4��bJ����^q�EZ)k��軳��5Z�Ŭz�Jht�0kqݨ�w�Ǣ�y+������P�E�P�Խ����	'�!5���=r�9IX2��&�[�i�["a�{]�ӧ��"�ꟿ���+R��A[޷�6:�J�D�4v7��>�5(3�q�D��]�3@f3gY*x"ڢ������e9Q��D��G�2rf���e��o�9��]��e���5�y�[]��rtY8��&�.����X7d:�KoZ�@Z�q?��1C9�)	hc� Hh������@7TM�R�m_U�ցL����I�|y�$oZ��&�du����4�/NϟM�i����B�/p"��88��1��.����ߔ8���,!� ;��Q�<e�����v����ړ?��>b�� �k��θC�'�~w�������4�Q��Dt�����j��*֙q��x�Ms���꺶U�ώ�k��n&b �²�=>�ٮ(	�Y����eV1�Ui�.��3� �9I��D���Dʍ�̦�	��������s�&���,&�UL��*S�D��Ƃ�����kBb%��s5}��Ԝx;�����$��̧h�~J�D�[ ���y�]]{s"�6c,�����:�G�3i���Y�q�����`��F��T&Ҧ�����K�L�M \/�p�BS�q)�&��[�go��D�F FO�S<�h#�eR��Ki�;��Z�2�%���J�Ԛ�R��Y��V<P��H4Ƴ�Q_^@N\�k�����~�dh�1�~�C�����MO>���p�3�����L��g�Q'�"+D~c�7+�i�u�0D{y=�/ �Mw�!Z��|p�b�r�|@����8Ī�����+�"A
���^W�"Q���:���?��KZr����;�,a�N,���掍��yH69҄��O��o~�7qy(1zko[�#~�;��$,��d�2��4�x�<dƟ�]%���a?̟'q�^�0�,�Q��x"�[gvu�651��xt�ӊ����wH,0���F�
H`��Q��|j:>��Z��^��@x���6B��L@s���mQ|L���(T�6þ��^4	{��2�^�^R.�pY�V��P!��O;�(��+�2��G������1o)���"X�s�^���F��䟺���w�c����Q����G�����*��. �`�}�&�xoW���.�@��1�h$�R(v ������NR���l(���E �{u;�W�I�n+QZ�E�J^�N���[�R��7~v%�.���zE�م�+�wO��^�8`3���C��K�Ҧ/�k���2�䣪��TF̔���@ۃ���6�������(k6�J3nc�����Gn�{��5:e#�������耘w��ˑ``o���2H[��n�Eb>ZT�g����j�]�tV��
J��]ĔP~Ǯ2L�\u��x͉��c��U�^$��$^ʅ>B9Yҵs*�?��:ƕ/2ax�3�{�^fw�(\h�U��r��d���A�꬧�Y0I�B�Q�]Z��E�y�F)@ӄh0��wL�9��9h�FK�?�!�)#`0����$��S���H8��O���"��j��醕�1�����	m�vsFX��8�.�N��i��f�,��x��dǫ�� �ã�r?���i���YYc�A�p.�*;}`��SEɨLbQ�ȱ�gm��]�����ʲ��?�k��#Р���*�,��C��;�АS�ƚI��vs�#��8�L1rjc��\ڛ����v��C3����L�Mx�'7�F��7C`�rf�LCǦР�=�no���v�V������{NȿRԟ�R���cI�,F#k�w.Y}<rIO1�W�kS��"Fak(��Mާ4c��t�p�=d$�p*ٽU�Ú���&-T"��p�<�{�=0���~B²f�)E��2㮀
@@iIu���� ,oPu~�q�h�j�&b�$ER�����J�S��H��-� e�T�䂪L����O�Q��D�]㎏�)r��IM*���b~H���+�u!�;q��%^n��M���X?Q�ܣs��|�캽��F�GCJ�v)8䎬�B���R�'�������'/r�L� ���`y���xM#z�s/X�;{7Ӛ����b�{/���I�硌����o�}�K��w[E1��!}:�-���9AD+n�J��3��G�Q�A6&w��*���U��w1�|N�D:���Pl`H/��<œ����5�ch�])�0p�:�+k���d��������r󑉄�H
��Y8��^d-ڈS���'���s�;�z�m��5�n����y�#"�n�ڗmO�#��,���`eV̔���v�d����[ �TNj.�o�
O��,g�+��Ƹ��k�J퐒E4�s�}$f����V�VHT|��Jv�#�}�E�%)ނ��)�砗�,��	���$$�M�.v4s=m��3�a�ᢱ�ERl3.DP,���k��6/n��p�N���F�F���d�	/�G��}�]��I������!+ o�]I3y��a1�;H����]		�S.��xT�@���[�G�'KI(j�f�hq�w�