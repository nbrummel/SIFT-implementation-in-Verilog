XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���P�2��e#���~���K�PWPX`'ۊ����B �!�F`��Θm��ܩpƐv Cn��N]TO�EɼA�W�w�����y�9/
�Cg�퐳*��aQw�7�ڠdզ�5ܔ;����z6�q��$?Be64��e)8�H�Q8�!�N�!ǌ��ן��JQ(;@�<4�d�S�� 1�3��y�K�Ѻ^�7#@��2Eࠚ�ɓ׊/&�8�@T��S �8�q��H���g��(������~=���}@��25�s*H12{�_
9J<v�E�(���܄�Q~�����	�H�t �;A��i>u�<��Zy�	t�k��H9$�.�X��q(-�ߡn����	�Q��o�wy��;38KmK��o�AoȀ�s9�2��׈!9��F�̚���:�b1�8;,!\M�d��YozYr<2�L��5=;]�Z�4A2*���x=o>���A�!�b�ؓ7�Q�����j���;9�2�<���/
��qnq�4�aJ!d«��*}=)	-�^&�"i��X����~;Q�{�Yg+���}���55�P�)1�q����Uq��M��U����3����Cr�������|�:�h�E�U?���6S6�TUHh-��kr�<���Ƀ0��,Kt��^�c�D�j��Ǡx�6��FP�D�6|i������8T��2 ƅ('8�s�)'���BpXM@v�e��o�
ݽ��HL1u��NN����&�W�� "00O�'�k�LP���9	d����KL�E�XlxVHYEB    15c9     850�u|���>��4IωW�h���XS�������rcd~A��sȟ�ۧ�ֆ�<-���8�����o��myߛw|�-�[8�GJ2�xרs�S��A[�c��R���r.��|�2<4���-'5��Y��0�&�d��=�)���}W#��V�{�t�r�?ᖸ��O�W-6w{ʇ��@��˞1=�B� q��[���������������9��ɏ=|�(}���**��C�Y�~WoL�8:�0בA��G�?�b�hZJc��2���

U���N��ʟm%�V��C��h=BR�rX�v�������x���"�����	&�!��ϓ2F����fV(�E<��J]�0��������훃��'�h#���plN�$)�0�$!MZ��}7򓈈��Mp�Bg�� ���f&ڬ�����r�4�NCR�/�UX����B�R'�B�D!��;�����-�CW�
9F�)�ma����d�������\<\-����%�@�P���R�c��be�����h��
���h��
���3�ߩ�01P����q�*(�>�_���k�J'��=r��Ҁ;ϭ��V�(�R;ᶙ��d�=��"���ƅ1��u�o[�{)���GWbk}���̭��V�|9� �<=ӓP1;e ��3x�uw*x!�ꬬ���h�W�Y�b�6�<�:� �<�#�����E��G�=�Y�?;A �_W���	z���u���lfU �wV�D$�~ԝ(��� �w�(�}0.�-��Bw4�I�j�ᨲ���N�d2��'[&0G�Y9U>���#d�7/�@�$Q�_�����k,&�9<f6�3ٲF�ֈ��i������vi�k��m��%�µk���̀�d�ޗ���a�-F��x��$(0�v.޷)a�
��Ol������'�^JA��] ��w!ݾ�Pd�ßޡ�u�;�n�qA��f_j b���P;��_�����cu���X��h��t��m���A��qČD���.:�]�㜞��x��t'�Kc�M=z1Uq]�m���M��l݁��m	-(�s9ҙ�Nܙ]�~�m'�0���d�}�)K��җN��+�j��������<M���c���WE�P�/��e����v�<J]��'�Q��7S�$i�˾ƕ���=Vr��*T�"�ĳ_-���s
�2:po�@[��
'Hj���*�#�
2�b�ه�a�P�i��1^�����h�_�ȃg�3���6/ZsK�u��`G��#K&�9��v����-�K�
A�C1s@P��Rm�\� �"j.��'(s{4���Uݒ�+W!)��)	��ě0�}�����!�6T�*(+������l��*�q���eҋ���L�����ʕ�/�7VsvNF]���`�����5��LG�z臷Tvgs��m��7'��'�/)s��秉9�-��׽|\�E��D�ThۭI	�c呇Ħ`��q&:v�x�z�T[\�y�=:m�F%�4/D����;�0N�H� ��}Y6NR���ك]��P�9�C]��5Vy�eM�����r>nӕ	W�����F��9��j�gv���閇������)��>�?.�T��O�ꉝ
�3+��CS!���N�3�'��yBt�}��ܝ&6����V���2��N�?d����&"c�_��>?�vg�/>���K��Ѻ2�wN��c~�O�-lv2��I1�耳>Z�IQ�A�*`��o�p�����9Ea��נ�
��T��Ejm��K"?H ����N(D$��HP{jskI,���E��r�0AiJk�L�W��V9)�(�	s|O[������R�_b��?ۋ�5'-�%s�o��D�J �����Eߩ�=.�ij�9�:o�JDr���II���O��Fn��0��9x*���1�9x"���d� ��e>���~�7�1r������!Wf|�>�X�w^
!V\�GS͊0�N�`1]��1E�g��p��-����ww�~Pd��!6��5輱���è����߅�R�Ku`�+��0�V����|Q�ɼE���!���5M�)�!*rF���D����$WGZaߠ=�a����Br