XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!R���9�1]��gP�H����@���1զQ���]�G���Fgw�+�P�<ak7r�-���n)gΑ�ɢ��t��|����5讐|���H,3�>H�V�jT�#JR\�-��/	��mիJz>ۇ��@�I�jڵ�	��K�q�?>�j�	Z��1�lB%�
���4G�G f��lq��/6�W(��B�=��b�:���x�`����|�?�Qg�6$����u�s����m�4#G
q�[	YX�;C*��t"~0����kЙ�h���s*V!���s`��Ƨ$h"�0<���������[����@/��� �Ϯ�@b�-/d0ԑ�T�mP6h��&!)�������Uz$�����q�c�k,�FM]EL�F�:��8�ԗ����i,�����<g�(<5J[p�`Ө��A�nl�~@���j��w��P�i�}pP�w�_�P7;i���*����@�T͖܍�ȍ���� SO1�R�oM3��w��2zw�tG+�.mBN�;%�,��6�c�����L�������H-��z�-<�
�a���N)���������z��A���#l����<4�xa6^01%I�T!�~�3��K�Ѽ��H�.�|���Rs����C��s�%��0~�����ϕ��W�jH�}���4DD�B�ۖ�ւ(��ǒ^%�K�_�)��Tf�Ǹu�`��%����F�r�I|��["������8�]���&w�},����!H�P
�b OXlxVHYEB    63ec    17e0Tc�׸�m�`��~��t�k6?2���}����e�ݤ(i��/�CL��t���}=�ֻ��n��0+�I�� ����,ag�ň�=����Nq�ˆ
���>�H{� ]���rK�#�K�Ͻ��b�n;˛��Tڱ8������9����ez��m����I�Ǧ�j�%�m��H�s���!k�-�|�H�}��Bq��Sf�B䳰��Y,e�!�O����m��Q��>�J2��{B{[�-��j�hq��K �oqn�#`��9a=8a�vf��\�g=�/ޘxM���f�w&*�jt�zկ�C��QҰ��<������A���D����&r �ɭ\���[�@�ş�&%(`7��Rs��7�Ͼ:B��b
�G���#��PysK�������F!P���1��XF��d�	.ODR��o�����1���󟕃�< :\d��Թ�j��-�=�ֻh��mX�hy��Z�K@�s�RweȚ�Y$h���4	4��l�H�r�<��08��7N9iH��65 �!������P�̪�[�_�.n�j}�Z�e{v< X&�e���S��.|�'ռ���5=��ݕ#mK�Y_���ͯ̈́Ŋk�E���a<آB��a��#���s�!�Z򍢔ľ�1���_�~�O�T}w�H�R�aj`�AߪՏ�Y� /���J�A��D� �c�b��YM�������o'xs�����[�x�pk�Фv64*(��恵�~�{��'��up�oڂ�(�S��ס��D�T���R1K�mh���[��׺x^M�o�t0�%o:�r��߁T�A�6&vp�k�{�)�?Z��h�P���C��
�oF�׿$�Vʽ�R�D�;�u6�������]�}���%qQ4}�T�y�,�&�n�T�� ��� �u[��n�1E�F���� ��0V����Zpy�����d<{���z'�?6��T6Nŝ]�0O���,�
�^�a}pY�v�/���7�����&L"�[x�G�I��)�v���ވ�r�^N�
�=�Z��DI��[��z��>c�b8����I��Eg��z��裕_@�mJ�a��M�x4��x3(є���~!TL'Zma��������RZ������`�RHK��#ⱟ�A{І��fyG��#.Q>N,H|�@lN��q?E�K� �������KJ���<��w� ��[	���-~zb�y"t�B�%MC�%�Nbo��eR�vN+��:��5�P"T����KX����d/��4�~���X�^�vM3���Z־d]IDԇ����5L��%\����Jm|��{`i	���S���F@�I�J9����`�`/�R�aE��y"A}`9�!ȇ;��Nte��z]��P[1���;~�*�m�R��5@E�r�A{��PJ�<ƅ�V���8<7�J����v���(w���k��OR�h���I��(L��vb��!�$���8��?6�O��-�X<"�
����z��z��	�����@H���Q��m��`����<L��5�~�i��ص��؃u��u��C-1�>I3P�$([�S�7R@U�q���/�S��R�GG��n�X���m��R��.��K]��r�`��݅����ƽq�X�@�J�غT�8{�ĩ-~s��t�ղ�0�Р\���Vc�4y����6�С%�vϞ��#
�ꪽ䫛��Q��]y?�N���Jx��H�8��Kvlq C���%�Kƛ���P�35�8���\fvP�}��Fy]`�65�U������)�F�2�ˊ d%r���U#Œ���R�MϒR�C�K��c���Y1�r��j���.�}0ԭ�?l.p��,�;�EC�Z �/��}��@�CCL��
w�~�~�\��o#����{�;����D*
R��p�`�{R��<:tM� =֌B��v��}�y�b=(N�	�y�GtI�m���[��#Aw��q�@MJ�2�Y�m�֟�<�p@�r�J�t	"J���ud)�QI��)�Л�>+��b��?7ks@$�(�������Y�-������Uv�q]��f�k'���K�yff��.�ϩ]�Wq��@�2]��eY����{�����C�%�Q��hR�D�dĖ<�����p#��s뉹w$?��v�`�����,�j�칹s@�a.jhw�<b�N���(Fm���P�2��3�&=ЩY��@!0�R�0�xX����_1]��)�y����,<������YZ������$`��zG��)���<th�$�U\��6�	^��:�=z����k�gUAZ�to�k��_��E�t3P�'�<5GI������G�&�[��r��$�:��s��(:��jp�ׂW�͌S{��M�Q��O)}�n|0N�FJق��?��x(R���ӕ�����������K��:�~�{� (��F8M�^W~���歃���`��1>��I��lv�.��pt׋H�0�Uږ�L9���^���g'Ǐ���3v**�+����c9-�Ӽ���1�Z��k��cf�=����$�'�	�$���FTn{~V?��m�b��_=���8����(s��qpcxG�Q�Hܡ�����g5Wv���ʭ��蹤�<���6��߲�_��t���zZ�B0��ȭ��R����}�J�X{Tdv���ڎ��P��|��N�,���;�E3e���+��/n״��j�-�'C.�^#;��<m��r6�D����O�M�Dq�hw�D�By=�K�[=p�/^
�l��ۻm��������=���1U�}��ϐ:R-1I2�����ROӌ�Tc�������w�*2��9��Gڔ�����cf´���L��]v��T�bdO6AQXEe.1,�^{�����o�9N��	pJ�k3�_���V�z�dV�6�.�ߍ!����<� ��j�bA���v2�Pi��|f'<d��&ꆩ�zO���S�j,��8�Y��a�0��r!����K�䥳��-����mk�=����bD��9d#喑:Cc��A���=f%d�	i0_Z��3҇�&D]sL��  ���֞�!���I�5��Jk�(���)���-���|�J�P�-@'�Fm=��цq�t�ki[���y:��Ru�5��E1R5�T���F~p��c���#5���y:\2�?Hx`U8KU/Y��j�C�j� � ����K�xN���`[�f� 0��%�ã�]G`HU�nlp���څ"ě�Z^���o�W*1�@��%���(>"��p���#m�t"�h�K����%?y�#ӟ�<����e�з�� ���F�Av�2��>`�B��L!�(0:�Q��Hql&�xө�h=��e���oU�#p��_�*uj�����h�[�/���X�nC�K��������Z��t��6���Z��sR�N��C�J�\J(��<�;b@#�e��=V$س�$�$�Zu���KM�/W$����-ԛ��
�XJ����;0n(5�Y-)d�T��[�;
�ub$j�`�L}�ங�/f�ݾyz~�-<�lΟe�?v��W����p2�D�;+c��K���0٠��t�Pm��(�Kl�(kw�Ag�DտG1�] �'EgP���J��)�(���^z?m�R]�zW4���Q���q_D�?�
U)���c��j{�i��8w:�t��23t�nG��Y�VY�΢�5(hW?�	c�����g�)�9��9ƟB��:�!:욆�Z��Đ5��e��L�6��|b?�E�_��G�~����������Ϡ� d��f���=@�A7�k�C3��)7��?���[�/��%��{R����+�Q��B���+���� b��v���t�N^�?ڮ%���t�w���P��ǝ���j[�

+��HoS�~q0�#׹�o�Q�+������ï�J�#|��C^垼?S�~��1P$b&��*�(���!{Rq�7����;S�� �%h��4�'�l�#A���]��R�s]�>���	�"`�����_�=@��BA��_�a�aw����Y�3w��Z�+���WxR�"�Ħ9�T���_���^2�����9բ�7���Ƽ�G�b�jn��'�o�p�e���ʔ)}B%JC���*����Ɠ������?(Wљ� �>���0 ����޳�PɎT���R7$#��~B��*+���!��N�el�V�83�/�� �>���l�뜏�@u�Ռ��
|$����Ʀ���5��\�%//�}�ٺ��+z����@@�jˇ&'Obzf��i�(���ۡ�I��Q��fpCL�7>�JjV������`���kb�S����֔����MG��̀�ʂ9<9��$֚���L�+T�����#+��#W���ؾ��ކ �
�r���#H㿡�a2�Jv�'u���A�1:�Gwԩz�LWmW+8UߨO թd��kf�5���@]< �D��	nt��}�%�P��� 9�a���.��M-�R�)B:],/�g� ˻A���u�"@�}k�����Ɣ�0!�S&��P-O�Àk��owu�d���̃�f�j8�.�;SXH0E@��ޔ�xa2)�C`���y�����>����G�7b���&�݃O/Nvy�M9�n0��$��p\����_J,J�:�V�-Bj�Ǵ�կ���#����d͵T�3�^;��ne%�0L&���K%v �g��� /�m��M�De�>�*pP#�6��«N���9�A�4k��Ü���i�W��
o�䦳hH�Uq���j�Xɽ����A�N:�@=?U��d�%#�`���p��D��X�>j�����
�A�5��3��bC�o.�d�?+(+�2���}�El�� �v�(�mk\��*���漢t\*��6��ک_.+˪̺����G�8��S(��A��"X��V�G���H	uX/.��1��ނ�)gs�[�_RfiÇ.����|\c<GA�F��y	0lT��q�>���p2� Jp<'$7��,�H+<ƚwN�oԌ@%B&�>��2$$���C������f�YE1Uv#�z9j��U5��'_9f��B	�*�͖
� �W�����5��kA�B��K2�8� �S&˔��4�q���*�=q�E����`H�zx�Z� �(��O�)���-�0#=.��;F#�?�q�ob޲��N���2���-dsǛ����N��� r9�t��!G�~"<Qd��ǙB�o�X'��NB�Ga��y�$�U$@�[">�y����~z_8;�{l3�Bw�x�x�&<�|�O�P���ɐ���9��/G�ާO)�n�.P���5�a�v������aʸ=mٍG428[R9�>߮�8�5�Vf];Mw�^m+������ћ�N�3#��:@쭏�Srkq��n��b������>$�!�Z��s��S1��3�C g˸�U
�^��^��Wdjv������+�#���oz�N\�7V�����s�V��HdQ�[���]��;`V0g��BQ�������,����)sh�R����!��:�����c�zws5�M���^�b���6w��� \�aR�{8ٹ*T���p�U��s��kj ��a�>
\�]�9r�$�!�@bC�Sf�׹�[���g�짝�?�a�`�����7�w{C��kHWg}�Mv�V�;�(1���� Fr5b������><�y�9TP�$��F�־�{�Z³�ݼ,�A)��;�S�rH�inXV
�e47a���&�~0AA����c>���9c6��RQ�� C��'u�l�
�E7�7��Ü���o��ϙ��[�e�!����{lf��#L�.F�'W�.��C�3s��ލ�� �%�������⊛"���V�8�&����좃K��F��>."K�\n��7V�Ά��a�K�����eS�	E4|��7���$�gئ�9�h�\�q۝U�C�a�7,�gH����1M��N�&����
�O\eF)�P��ŵF<��dL���Y��7�gma�m�HA�^d�Bұ6����������f�_