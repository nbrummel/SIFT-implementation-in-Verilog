XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i�t� wi��.�X)��m�h�ee��9��q�aG��6zb�B JUY����N�f؇8��+qwq�8b�g��њ8~8ዬ`R��{�*k�ج�[�kʉ,��iF��)@fG�'�4fd7]~���0�e�9�h����'���rk�[�e��:�OR�k@��z� ��6�z`�P�8K$�V�&����X�6�BZuC�K��=q���C��2Ac�uI[
�I��>�L-Bt���C$����k�?������P%�e��2���{i���j�Ra+�b�<����ۂ�fB"Q����]�W(iV��a+�03/8�N�'��sQ���{�j��_X���	e�t̑3�@��>��>�����1�-ۮM�]�W��uQ_��l*�+�y>��7�eX��N��O��0Y��&�H�(����d�^8��x.���z�^n�꬘��Z͜n�����vq�6,�Q�75}Z6?j�8� >�^�;�u��>���`�-�Y��-��J7�X�w�a�O饤Y	�r�؞3S�s����.h������+��Nҗ?;��1�F���[ɾ�
�����;Q#�H9=�ڊ6�$wP�o�S�N�'��#j�n�&�9*��1��g�ĕ�A�M�S��: ��^�-�3>�%�_g��"]ot���ˉ|��ȠL|:ᓧ^7�����L��jD��{���K�!���xa:0X�9Y��޾3x��������$X(o�O�9RJ���=wR�Ά�K3�XlxVHYEB    b8a6    1ac0��X��8�f��4�e���	P�oHy�ƴ���d�6d��}e�l��!<��ex�WL�] V��1r:�IHh[h�7� ��)Y���V��n�G"�ߡ�ޕ
v�v#q`!�B1���͜\�W�ZeP5�zA�� .������(I��y�c��4�$id����ġ��Nj�%��1Y��,�Y�9�Ԅ8P�zʹ��JF��˕e�^Ȝ�EX,�yW��wq�0a-klrgD�M�"���2�gw��j4���f�4�Йo8�P�.�����_S(�~�wV�xUQj�ONL�`�К<:K�> f	6���ä��
n��~�����^�-��|���k�1�Lø�a<[����=�vy�ͼד�ZE�]�]]!�*j�_u�S���?�ln�'�<[�r��LD(�xj�\���kB��{����f2|N���U)|�B������X8o�W�\�	�#�f��0����">&#��푎m�#P��ǽ'�o��6��3S�OG�pH�5��$�$v_�bE���&F_Y+e����\
ي���?u�D�Z"��S,����%��H��!��I��i̯PuT�&�9�0����~�^�d�Cu0K�xfV�d{&�5��m��i��<q�ǖ,�!ؖ��(���p^�u��X�mq:O���������'k����g�w>�:�2c���!\���P�9����--%�o�3'zΖ��y��X^$=Ӿ�ޠ�@G���v�OwP�,#Mj$��hz&���Ǽ�� �+J�C�ȒBEXkA���} Q������N�^��V��3AD7w0�#|�������O�8��ʆS�k�o�v�>2��D��&�W+���gyJ�Y	��o���d�lP'��q0 ��=��*�g�y��\��E?/`E냜�|&!�NR��z�*��̘�s�� �gv9яh	q�Peӻ7(����&@�� d���WCtU�2~X�cX�
��z$Y�s��M֟��E>��XT�!��
a�}��A�V�bn sڝӮ��L��O��B�쩉qoY������֋_�	`6��9�N����L̓�
,?
���$t���K���0����oNE nX���:�d�2��O�����,��0�weE�b1\˦v՚r˨�����XN�&�۩����s�\������L�<��K�~��=`�?|3�ֻџJk�F˶�p&`��+��)N�a>�����"�\�,�D�(��4=��l�t���v�e���
��޺�|��� x4���?8d��?��ʞ�ڋ��`��`�#��'2G!����8�/Ō�h'+0�Ҙ�sCʘ��ȓ��d<)����GQ:�A�q����G�=��׬f�����6q?�[�<AK��?a��&>v�k�m�\ ��Ժ��?���֑K�h2V�	���=��M̈ᧁ�X@h�4���v�Rx������e���4=)'�V����b��`�t�s�+���m�r$c�C��?��2'�Dq���,�ۊ��E� U��.�^J�=�
췔���p�<�/���<����9�X�N�>�����E`��g��cb�t*�ΝnT���z�l���g����g�@M�<[e?é�i��g�/���nȟ�d�X���)r=����`A	��
A�.8jGĎ�QO��s�˵SKto�΋�K�ps̛�mf:�ܲ����ܦ�)"�L�d��(&�"��PE�o�nct�{�����Zv���ԭ���#!�����^����@\Љ0�n�9R
��M*����)y���6���#/ݻ�1�H���1]��������$�G�D�tZX8�����L��򽺖��pdj���7�(~��]�U��3M��� P�\����T�	[X���*`M��p�����us���>���r0?�^����6u�xp�H�4;�4�̯@g6v��_� *�]���V����ݣ��t��Ih]����o�g?W:>|0tu��^V�� �{��b�����h������, l��,O0+�a0�������(t�[^|^�o�h%ln�����d~p�Xup�	�6���E��G��j�)�]�q�ے��\Au+��OXkv�$�S�����;�5��u�m��7B<h���"�;A�cO(}�װg)��p;�}ո��h�K�>��_i�[�K�R��n����i��aD��|HZYd���RFx�⌴ڶ�s�&t����jU�>��	�$�I�nl|�Y��"g���������Ӊ�P��0/;C����z+���)��W"��C�]���âL�&���G����t�c�ִ�#�|ۼY�AIV��!��cr'���zǙ���p)}�ٕ+�9�#�l���{�]un�vQU��%�Soo{LIEE��(і1�fnm��W�w5��L�.�V�<�c$��[�P��DC���-�s�:({�?�y�.Hn;�GgD�nL~�ʩ�L��S��!�!MO��퐼윈]$�v�0���P�5�C��	�����n��j�-��d���U���x��*����u���eQݛ��aD ���r�6���ѡ�XV������i[�R\�gk#:'x:f�~G�/SĴX�|'ơOԈ-���.���agb��.��h�;��H���(@7f�R��RQ�ﾄ%?��������CI�`A�N��h��ѡ&v�W\#�=�Ev��|e˖�[07�mg�IK���K��]gxl�0���V��ģjZ��lk�Bl�4���y��|�X��X!bHuG~�4��n�$�M&�_�����!� 
����Ka��D�
\����asΛ��aP�w�
�5�bp��w~��ZF�Jvm܉�^5�	����x��|E
[];4�t�X��p�!A�jTw�����P�>%9��ύF+�G��[��9�e��R���<�{�b��u�����MML�2ʄ=�U:�L��s�^�#Tv�1�gI'eѳV�A�SJR���7\/��u�f��>��W�LB"Q��{!˨T��!��^��"t��'^Yc{�a��OtՆW�����%���Z]���~����&{Pׅ 0�"מ�Y�jVb�XY�_��.4�s�{hӱ��l�Q�	jj��0� <ׇnK�%��tq��D��I^�g9ģ9��3J�@L�|M��R{~7�ݡ�E���D�����k�a=�y*����ݕy��&B�r������H0��e�[,�A����WYY�#d���D�Y�%RC+�͇�ݦ�?
6]ϴ`����h���<���������._��� zˈ�r�80[���]tϏ4!���iG�����s����Hun#U�ΖU�ĥo���24(��F���<����7�n]/F��1�N�@_͝�|�y�ա1�5�9�)�!�[���'"\;�X�k�\v��K�c�Ǯ�mA� F�f&ێ*	Xy+^�����g�Ϻ�i��9��N��)�X8tk�̐���Ʃ,\���icE�n����R@V\1{�qtn���TdTͅ"y_b
\r>���{�^B��X�g4�Bk7�熨���~��AB]�QE�WL�C�q{G�;�B�1 �k19+�1Fв�>���N̔�F��C���Xbc����i.%	��J���I�?�l��G(�)R���0\S��c<�~A@� ��}�!U|z�;��k�EoYo���e��C�?, �2,�S+R��:(���q̗�jIO��H�po�g�65�2+����9<ʉ��(�8��8v��^:�l�FO�a�j>;���1����eBR���6c�ML�b��,���n�LU����q/�-�1�'��i��r�΢�U�j#�t��/�u
oG�e��*$m6t����a.Y����78I(�(�����ȟ���y��Q�{.���c�;tM�
�5o���h�Z����ʮh������?o�M=��3ެ���^'
KY�I���:�\��b�U�Z���*
ջw��7�b�g()	�
-��G%���B���"�� 븕I�����}B��f��1�&��þ��}7U�k�����H�+�H�lxƖ2br��fNۀ0 8ew4��`�Q��W��ҿl������f�N�q0e$(Qũ�#"����cD��&� .�V�:�o��_��o՝E����f"v!L�Ժ�n,�=�߳;�U����5L6N�E)'@l[���b�v�5U�,�f�� Ex-, �+�/��K�LL���	���9u]�JPb@���o'��._4>|i�FOGQU֋AC�
h�%2Hg�N�B��o[Q{5`9N.`�ӝc�3�V��Xݶ�3�p�J�7��uX�nC@��MS-�G������!�SO��MCY�JB�9@U��ms~��U���M��]�:x⩥ah�Ħ�����L���m:�v��m�qC�A�ON ��B'��N��p�m�l�-c�SI��>n��G.gwsH���������a��F�8���xb��3'g��8�OU��B.��2#���.�\i�����x|�vY,D#�d-�n%���Ʉ�fV�t�:E�Є-��E�S�|��е��CO4�\�iA��(�Qk�{8��w.[.G$�E��r��xӬ��^�G�e���D�Ǜ�*�﬙P���l���f6��T��r;$���/d�hs�vFH�JeY"^6��{�8z|���`�ԜuڬB����X�b �l�̓�u��@�H�!�)��T��f��E��ҩ�������8���V����OE���(=
�<'O��m60u���J��+y���1<>ѾZ����ĐP�s���Te�ۇ��O )��ZnP�$JJ��l2rW/"E	�:����9�Q6��a�Q��S����b�]K�=�Ē	��֫F	�10�߼�!��T���\�J�ul�[/�z�G�q��a��^�6�Y��[G����YtGa���X�m���I�����H�_F��6��sr rylG-?ul"6w!�G�'I�nˠ�i{�(++<�Ҥ���%�D)>l��|��ǲfgOͬ3�OW{�!���!A�;T������/P�t�~ő�b���k�&�[��j�",k${���m(7�諀P�ґ�>�x�\&�$}��M�n]dO�s��V�'�]��:�	Z�j�ߐ+�4tש{�(��1��$��]/H�/��K�!�N|��GX����H�j�e�C���۫�4��xMg�e6��M/i>
W���Q��-�
�Uu�ԢJ�<m
�}G��`��[�Zչ���E;�H�\R�pc?�b�ޓ���	o��7������-�iz��ڏ�p��\�f��n��~�����k͍K��;��r�H���:��`�����z��?�k���AJvt�����K]����o�X�`���S�wʿpg	T�Ol�F�?a
lC��Z�n��T_8d������DԄ�\�""DӸ��K<�|߼K#��f���es�?��޽d!��i9�'\�̍�\A�KҟҠ��mĘ�*�!��������k��@!�ػ��gs��S�~h��j,�وvĭ��_l��U��b|��A:f��z%��g�+���!�����-6�n���p�rE�WvN����\��뾡>}�d��v~2Ͳ����B�k���D��a3MڤP/r��R`��	�H%��@�2����S.}�ȮѨ)9�]�E�l�BjD��{�ދ��f�p��%hDj�\χ:1�T�Am��2��+i��*k�S̟�H��Ҭ���s�,��?�4&9�ErK�s.�Y��;��8|��5I\��Q���2d�#w�}9
L�l�uz��7�܇�����mUC���kScB�ML����}��ò��W��x-ĩ�@M�!#|՘����\��x!B����J
%�f�P��|ۊ��G�|��}�C�o�n�2T-
h��~L�UX�P���)���*4Շ�@�e��u���pǳ�.�#�e\�}�c�����7�9��.K�I�[	4)Pz�ZZ�{�� ݀`����
Hn���ՙcv���b�<�q��@���x���L�#Sl>׆�;j����a�*S�|$�ӝt��&���;g�'U���8�:F�������\s��Z��i���pry4]��L}�8�
L�ϧ�`=U��T�Z��,N��0}TgH��4��#��+ʹ��!K����B�=E�AwF*-���� ���;�K2�9v5Ƈ�����D����=��M*0 ,R��죑*�0��7�h�b/xT���\Dޖ���!�2�bV�����jξk�L`f�?�v��v��t��k��G��gb	�W�L�p���0�O�*��^��e1β�	Z�D]����g;׷h���AM���Fh��d"���:��%e���;9q���;�t��n�R�o�`2#i߿
��:h��RE<>�ԓ�3�*�x�4���MjP�TO��ݐ��d@�q�W�tcA� �ȯTÍUx�ᄨ���bA���1�!�P5b�t�@q�b�٩��e���9��o$�f�Q$���'�Iq�d�ڬ�H�7���A�C�pX���$�T.�aS��"'�]�y�5�"%��:t��#��yӷM�Ɇ
a�WQ7�g�o�|��ꨲ���EptU�6�/F��>�3�Ex�<c���*���НI��湌z��)���*����Ot��TPMb_Tov���oZ:���O�"���Nɩ��P��Z1���5