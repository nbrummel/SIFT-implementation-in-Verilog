XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t�������'�v/�0��6GXh���S��"�T5)���F�N����M�c �M],^jܐ��b�WC2`����Y:l����S��L?�s>���<&�Ңb�<���$$9'l��;������jXzT��j��$Do����\hU3�~e��'u�F�^j���BӔ_��=�Z:$��
Ф\f��E��g�Pd�oT���O/!Ų���������b��l}� ��q�����H=�Hn���)�u�ϱ�ރ(��KV
t{�9E��\��G�S:j.͑
�h�Kt��K��D8Y����t��O5�=�nf$/V�F�%����0��h�J��%�?j>�ފ�f���Rpe$K��erJe��p���]#����o�֣�x�`v#%���/����� ��O1����N7�������ga��w��������,�6,C��8�V]U��INbckm5,+;�~����<�}�+x(�������5�͖�u�r��;�52�W̓r|���D�I{\�)Q�c l�������E�/�	��17R�&%�����Y��7;�#"��#����P�-X��L.�l�F��@�4�L���"�@�����S��#��^+��a�4S�Z��ma��f����ZI�:�4��XＴ���X����-p�����q�k�� �g��D��Vi�t �O,�U[cr�:����D.#���O�3H�ږ0 *�	R�
��UE���uv�d���],�����TRu&|��XlxVHYEB    549f    1060�
�9�^ߔ��U�ด��g��9�(��d�:.g{1v�d#�P��*���iIr�eNP��Ft�C��p�`��xk��H��Er�p����{*M2����At���WT�ٯ����'œ�4� �3X^���~H��[��[���~�	ewV����[�"`4��9V{�#h�M�c�+h��;s�d�d�z�9$ԩ+��#�n�Q>�J�������n~��*�ā{l��ޝ&�ù�e��/�#�&;��/��T?���۩T���&E�A�jͯ������U1Dy}_r�ܴO�I�k_��q�DB͓)oAE6���j�ߟff�2^z�5�3�J���0�x}gz�,����a�����C�0��NP��~���A��^7	0��UryU��(�������{��(w0����E�ui�#�V�?@���)�ݓJ\Z�RS�ˢ�ǥ�(�%U_��	�h,	��4��T�@�߸n���]P$���kk���;���2)��y���OrUxbS��Ӗ�R�i���k�t��u���{����e�3��h�D^���E�?��2xVM��0�!Y��П1���1��R��G�D�޻I�XU��yL�x	��I��;>�7���6�|B(��>4<%и5�"�&.�(��/���B5�"��!l�\�t�:@wc��J+��)��sU�.K���ؙ`�!J=r���F����9�*�3Y�t�����<�[ӛ�x�zrĴ����D�6��Y�6�w��{��m����H>sh�QZHH�k��c��H��F9)xM!���cp���"J{H<�v���;@b=8����vq�v7�UF_KB��ܩ*�]�"	'Ν���c�O������I/�G/�^^k�s] �8���v�0^m�y��4���9���3��n���13��-� Y(���,����iʚ��@��RJ�+�>�2]s��������$�~'�|��i(r��K��kU���go��|Ĥ�x�~�. �G<���~�O��(�gg����D}�����9�eOL�c�D��$��o�S$�p�u�V�z��*RF �V6��p�y�r���^�-�SY�n��͐����7Q-p�K\4����/��<�"�
���@��{`�)	ı��%���/��s���̠y��=�;��L���5ZQ.�8��Zo���/���6�#�/Y,�p��=���TS9ԍ�ջ�Z_�,$$ �YT�2��/� v"i[4�ڌ�~���[��Q�-�.QG:Y������P��L)�h�3Z��>86"d�|��֤nx�Ǹ3�3�����.K�5�R{j��XN��� �Zv��+� !�S�A|%�"�2��k�R4uY<�	��]��*�5���}�w ��Z�&����[/}f���$
�&s�~Q��Q�L0�.2�mض���b�s�)A����П�վ(P��dm��d����
���ل�?tٔ �=��P0;��)�B��K��r����W�\�G*�}���^��H:zY���{|#C����g�}�JZ���Eo7��Z<X��g���XU{��hu1��b!,�Mb8�̓�� F�C$�.��<�V�Yh�@]�N.1�Q)+�A�i��|��B0�����	
,���c����7�� 	v��m7�npq�.�b�y0LX�V^ԝؐ,.��I�`C����N.��y��"�o��x��L��ΝU�����?:U��h�4���+�����mFD�hJ`/��C|2xv�|�9�+�e���\�C QzEWζg؇�	�(Ǚ�sao��2'/�q��px���1�j"���O���F��|��k�+���_��p�`��-���p_���cj��e�����B�^wZzi�3	��!��-��TB,]ᳮQ(A�P+Ć�7���oA��b-7k�1t'u��t�z7kf��#���Y�Q��§��D��gj%	|�Y����%]��-���#�1�-qn�(TF�G�y��Tޒ`����2���vn�a�j�����{̼쒁��n�==~l�H��O �Z�I2�;��1�4� �55e�"�%��F���'le�D��&g����QI%w%�`Q][���{��W��Yk�p_��|j>�ɨA��7��L�U`B���]�j?9��e�~�"Th��S6ʑ�G�Ԭ���r������J멄[�Iq ��Xك!%��ߝ����#;�"�Q��5�ݑ�c����OK|c��[��i/���H�"@@m� &
���/󝩳1�4R���[����Dy��.%a���m�Q���ыg@��M�;���"�[Mُ���%�j��Be���cw��2���7��6�|�i�D@*��Y���z��d���PVT :��k��:E@A��bW�{7:����QG��[��5H���ܻB���yi�<��,ꃭC&��i����~%��u��A84@��|�ν�t�Wb'�3�q�nx--0���q\�����D|�sÕ��A|b[�;��ʭ&�7@��Z�㸲ROb��T��Z��I�`@ �S�>�w¨^l�hIY�Y�t�r�@�5���!J��Ԫ�ny�����J���?�:��4ԏϕ*�וK�2&R>�K��T�y����D{"P�� �]��D+ak�3��)�M����JU�P \|-wZȮZփ�\!����el���T�Կ@���8'���Ю�8@�W�霘1���F����GqB�b�%!�f���g�����w� ���_�s'��|�-Ϻ
�E75K �H��d�	�.eib�YF�XxP7z]��H��=�L	�i<��0d�N���H����Y%i�)�׭�'�e'U|�|	�	�_�==$gZ��[`�$�YJ��tD�
Gt���;�sM��H�P_5�b)ǲbA�?��R�O��G�h!���c;���J� Ee���O[�%a��-��4�;R�s��S�1���HP�$9+l�T�5M��!!N~%��> �G����Ĭ��&I'��~��=\b�I���Y���{Y&��՚�t]Ȓi��i���E�b~O�B㛾>=7�f.9l�	AY�ѡ㣳TR�Dy4��J:� ^��ZPG�k��#y�[b��7��x���LF8g�#p��HlG�A�n���`D&�ͧ^���bQ�j萒���շ���� �)L�q5A�$]U��2�H��m#�ܿЈ��NR.���x1�f-�dD��������6T�C���G�/��I�����4���C��@4���(�矟N���N�A�<A`��h[<*^�o<���;���myT���ۺ�׭�>	��a,h���$rm�H�?�.���y�������kH�Ag^E�@�Kx,UDޤ��z;�ǧ��Ir�r9����7XY�pbg�������p3�z�炪�7o�Õ�Fp������#X����$��_zD3s�d�\���quu3���U�!!�b�2{ߴ�,����$bS�2F�<���>��)!-�2��]���a'm@Y�2��ny��n�����I���Q/�&����kޮ]e��c"���xJ�{��F¼�]~�ʶo�	.t\��ќh�`%�������م7,���5���&�����E����C�)��,U��ȟ,�o������@�6B
jAc0m�T8b++���{E]Y~S�h/�0�����@+Ʒ��rG���S��s�w��b�Φtdp0���Z�i *g5}��4xV4(-��vǅ��G�'B���{c��wV]�R웉_}ҟ�'i�L+��ԯ���?UJc�EQ\�Du���˔�*!���]�cҾ
C��LI8�&ߓ^W�J;� 5�*�e�y�g9��E�1O�3����p@�>?1�S�ҹ2aҌ�X�
�mf����Џ�@�}G�N�w��U6O��pK8�C���ǮX��h��CG4��p*"[���L�C�[Fؖ����U�4�y����Z\��@�����������QU�}Il�h�5��L�Z��H�p^�+�Z�[&z�6��	 b��V����|�#��b���I��r�pgdҒ�	A��L��D��J�h1�F�FS�.{v
`�t��2���&��3�~=�1�r���#]*팖�+�\���	���c���