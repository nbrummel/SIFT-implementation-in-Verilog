XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a���b�����d��p�0p7�P<z\�t�Q]��^��B�����C��F7E�"�M�����rov�V� ^ًȭ	[P�m�O|S��ئ3����:���A\m�q����y'�R��v�N�f��3Dv�� t�e`���C%i{~0 �&5��V:C���(��aPG�a�7Pj���Zc��g�p��lAUcdz�\a>\�P��ѹꧣJj4��O�F�z�w�L�ї0��~���֑BD"yr�����G�*V���7��`��֛�f�E_e���-���o��|*��ڨ���� �t܂�N�)�$%3�(�����G�Y6�H�7N�Þ|4@�w6�Dq�=6%:+=�?y	f���aZ7�9���H̫��&P�_a��D�duo������?:v�U 6h����0��*��Jln/@ەd�T��\7��6�bb�T��0�RB���������/��W�I����fX�p>p�՝�}V�+�a�eI�[���	�Ύ]��g�w�q���p8���;���kY���i˦.#ɤr|D��A ���E��w�\W;o�1ɀP���Ψ2�<P_�r�'=E���r���1�vPֈiV6yLx�t!�YR溇L=+*^*;V�x����X-:Q�xj�)J�&�?��G�(^"���l�M��
ߔzVһ/*�H�ͽe#Ov-�>;�������! �[�[ۋ#.����K���F|O>�a����%��u��k�V�ZT'�5��6U0u���D���Ho]K��`�҄�k��sXXlxVHYEB    2577     a70���q��p����qÇ���f�%�0pnr�`�*�$_�>��=1&QC��M`����Mfe��G²9�.��vZlѧs��s��R%C���v��XW��1�C7�S� ���9SC��4����vV�8���,�]�WkAsw��ʹ��2���oN�*_B��B'��a��ƴC��b���iK��T��vv,bB���Ye�KI��=SW�8'1���lW����IM��̜Y6��)@��� �rv��>��Y�sc*t�0�:z�������֧����6xe�4%1�Q�� �n��Nt__�{5Ó�^�jT��Y9���+��L��k���aw�+*�S�P�|"6�:�GC�X�h�8�ݺBv�����h���Z���,lNȳ���lyz^� yn]��~����0��^p�=�� Nsh�k� ��v���(\�6E�OQ�f�
��m����-,�f�$@8BN�,D;�q�;(ԠN�l��T����h���6l:�qW��
�9Y���_+����.1-�*�]/Δ���m���l�y���y�
�9���qc�B�>�Q�T�'�.߸�[��e�$���^�����#Ò�1����OZ�i&	aU��>������k��}(��H�OY��_�v7�X��z�pwR��KW���1'��{j�����)���Wު�?K��C�u�2�9@( �aRJ�5�v(���r��"���,~	�����y��z��Nnӎ�qC����Z���w�p�g�0&�0����p�?��R��oUx�l��}�iI��&,�W���R��C���� (0%�s��+�����l#y-�I�2l��������� �C��a��&�k�(�閅�~�9��C�N����y��.O辍�}��������KsW�Ż��3�x��4NGIE�9P6\T�#J���o�}���W��8�Έ��Y�9�Ɍ��(�,���͈L8Q�j��B��(Ǌ����m�-��}�&��O��q,&�����'���z�2��G9�=ݸ���2��,y���h����*�B���%Yⶰi���UoAX�!��� �G���o1aH�K"E�25z�Ľ�m%�͒�˾�� �]��b^�P�K:��O�<�o�k��=���AP�:('�?��)�^��m�_"���R����J��4��RSQ���G���Ƃ]���agm�U!ؗ1%����R���eq\���Qt�:�M1V.#��'�ZOt�:��\�x!��ZȂ�_�7&���hS*�'Ht��9o39��Iu���Xjg�jP�ߏ��Nꄌ�9Xà��"�f7j<�Q�?���	`꼎j�LU�t��d_�E��qoL��M�Ȟ�U�!/�&�as��8�A��p���Q�i�S�+�87�8�]<�T��'�܀�d����f��hE�+�]��wk���"�S-���L,h#��(��
wCx�^�!�r뾁Kx�I̕��$
������3�+��Ɨ��;��p�p�R��/~�"(�7X[�r�w�a<4�nD��R�Ĭ�
G��h�O���TR/'�-���1HK���T!d������"��1�{��[�,!)W�?4��u�r/��о���d�"i�̾��d׮�E���P8�@���B��~��4>J�w4"��. �x��Z|�	�{��R���b|�)(m����C|<���L:�Tr���@%|SD�K�<�������~J��Yk����D���pX��]z�P���g���y>�|�i��?'ՄD`����G���,�H 8Ox�:2�@�MT�7�X����+�W�@u���ԧ��z�w��t�g����	�0�%�Sx�p���%�~C��R���@��K������>����}��V��7	����čk���~�#��������� }f�ƒ�ƙ/H҃6�C�m+L��悔*SS;�����Xzd��q�ތ:�dz�("3y�Q�}�����&�;���ȾE�1Mˊ)���k���X�Ss[��wT�@�2����������5�|� [�6���dR���۬�������R
�����ҺE�,�)��A~�-Bb��7."}��&?Z��%�x=UA3~������g{�Z�{!v���@��W�p���5Y6`lM#p4�*�Q4o&U���`�b��t�o5hKsmġj����@��m������)����rx��w�����/�1��3},x�5��(��ϺѴ4����M�?��c	�R�k4��%[�N��3����ܠ:@ne4%��kl��[�bd�n!=]�	pV���ra��یI�	HE}��P��e�L�w����2���0�:�<��F��K/�G�S¬p@��OS?�8,�`�Pw���7��xH�'��i��pL����� 	�(�s�wS�֨�$��c��*i����y��|"�;�ҒQn֜G�A��>(�U6/�v���{K_6�W�
�A��+��{<^^~X�c_��I)�.��ޖ��Rdf`fh��"w&�|��*7:�9�
q�S�L���F�����G�s^��ں���3��q��# �
���!�f���)�c�t2���?��Q~�� ߌ�
�H�h�?_�
��_0�"W�