XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���L�F�� �bS��6ֻ�H��(J�d�J�,=`W�D�'b�W-hg���'�����d�mȺ�2�ą�����i�c��օn	��ziC?.7U}"BSPm���w�Y��ީ<&[��r�>`��0%"%��@�Gc�s�D>��	n� Ya�����]��׺A-�C����p�9��he>�C�P1�l7���<M�w���s0�ʌ����?1��0ԆY 8�Σ�0+��~P�K�%�i<닔�Ѳ�٪Cb��,o�I���/ʿTC��\���y@q�'��ܖ��o�#�f��ꡐ@��%%����`����z仛וB�$� �^z�(ţ�݌==��ۢ����Cఔ�A������CM,�
{���B� D������<��[PΓ�(]�g��V��h�;�����F1�p���F�@�{���h�V�@eP��'-����i�;��{���Jd+�V)m�M��"��	�&J"����WC�
�ǲKm��u-�o���I�w��́/6t7s��}@tfAzbp���{r��iB��|t3���U�v$���*�"Y��=��VO dԙKE�B�Vwz��	~����U����"2��_L�����{�ks��Ȁ�P
˲7��4K��╩/7_���Ʋ���f{����e;~��?��������2(�*��o�b6�W��k^N�����0�=(����A��f0��xO���!��t�ыqw%��l+��z( [G��[@0�꡹α��P:$f��XlxVHYEB    aa52    13d0M�LVGqڙ�C:4 `P5�G�� �S!HZ`�����V3����䁡�ax��W�R���[�U��g�g�q�֥Ax�<
�GP�[���몉+��Q�xi1X�	PE���8$��TqxN5ĳ��φ�ՐT�_Y.SywgA�ܨ��Tp��a(/��!F���Y|bv�����Ҝ����/�[� ��C��]�Fa-&�Ϧ��,�WUe[kp���c����X�g���˸�<FŪ$P���{�7�#K
cӺn���3�i��/,$��K!��ӯ��Y�~+�
@��k!TK��{�ٸ��!w��1@fn=+&��J������Q��M�
v�rj���Rμ�.�3S�{�l�g�,����υ��>ǧ�*��cw9�F褲��MZ��޹|��<~/H/���%=y��A~E����������%�U�en��)e�nT��7*�|����&;��a�������r��%��M���Ԕ���]�c&|�����ڻ�u/�Ŗ�̍[RH��^�U�w�ױog�����Ғ�ð��'�U:t�U�FgB��3�$�2����MUBmL8]@ň�l�[�D��50![�ʖ(��s:>xd�M�� ��1E��TzM�����N��V��5S�<��6�鏾Q��f_>���Q�뫃P�,wC�u��im��7H���x��>�O�0V�����QnLS�"�n����u���\�[�s��NMM��C�2b)�9K ����IL��#����i���=�2�=��<+�W��C��o��t|s��H��gq���F�����y렚QX� 8r�:�|֣�}�E��l~(b��Ti_ ���5��ۓ�z,Zez�1�`��s;�F<LNg�S����a�\o8�U�g�/�f���v����B@��6��O��`�jB��9�6]��umBt���H�����Kr����x��Xs&Om�Q;��~�y��v�pG#���*��K��1�ws�%S�͓̞؏)��/͗�' i���9�"I3�m.�o�1-�N2W8sc��$�p���iy]�0�7�p�S,G���9�ַ�I|�0�ں�HSݼ����۟(��Qi��`ry�����'�4a�M��1��!72	R\�Q�rk�n�q��'J����SV6��'�Q��N�N�Bl(Ǜ��l���}(L����Ȕ��S�
�v "�3�C�Ӱr����Y:����������Kc��A����n�lS�s��W�Qh��U{��q�������s~�b�O�0�ɝ{}�eL�' ��련|�ZO�0���$m���ޫ_�U���V�t�#.9-��&K��kl�·O��g7Z��4��:^Ek�ğ3��tK#����O��zj��v x���B��)�rd����D(��;���I��M������mQ�)l���f� ۶+p�K�9c��]����Zu�DH��rl��w� ���A8(��������7�9+6�IJ�fo����Cf�f�O��s"�<���).W<1�-�z4*�~48ah���!U��c�<n2�/��qh ���4��}�<+K�B�e�W�$��W��b)�W1�F��}�+��K��Ő�����g7�o��P��vo�6����V.W�oͭ9��ޛ��M��g�{��,Hɺ�q ��a~լS���Gq2��bwX�-��1�'�,���2�_c���I	�v�1�ڡi�P�x{_\�a�%k��k�����I@`(-ݧpE�J������*�[�B-�A���H��Q�����>���zA��֙�p�r߁������}��Ƨ�AW�FƮ�����,~ a4��w����V2�������`4r��
��t�<�8`&���q�B}� i|���1�R��������5�$0o��3F`}���o���k/ [��|��ا�c��M�9��G�P�B�ߊ�j������������9���*�K���jvږԕ��	�+Q�/`�5���ᢹ�@q��R�SVLx2��(��Đ=9-�1(QhP�%���C�lѩCZ�jy���O�)���@� e�ɴҭIn\�l���۷�f�",ÈQH�.�v�Ծ�w{�K��e�yk��j.�nXE���y7�ū��_p��҄$#H������ Iݔ�?�V��"��=#�V���z��%���+�to��m�d�V�|b��a҄ڑ�j��Q�-��Psv�Ԫ4��ۛ�*@u��_��Q'9N��J�4������S���e)q��(���G�T����%JϯP�_�u+L�Ar��5��%���\����f�ʤ�,���Ke!��\�b�� ��.6�x�18���?B4]��t島����U�\)�Њ�Y�U��D��h 0�����V,�V�Hv.�7�5�J~����'�@2��V�&e+��G��c�E;�%�mk�v"��k?z��~Kq�lZ}:f�҆p�u`���xY{E�@�`���A@�
(��͎^w6�>mdƷ�ev�c|�閍3F�B���h&y6�Ǩ���_��|}�
y'�����&�gm��uq��X��PQ0^]#��"�'�~{��X�0�'�`��Q#�p݂��,�&��� m�A�%É�8h?2#�� 4wъ��yq����-H%�>u�;F���x�1��ڊ7�~��&E��a�f�A�1i ���o_�	:=:����i�Gk��뫆���*܌܄�OҴ.�λ�X����nZ7��6_z�T�����#@[�M0�]��ֱqӛ�H�1�8;h�����w�H�OAh�V��5���k��w�@axp��h�g�>�DCI`�f%s�T�����Ы�,�7�V�[���/�c=�_��K��ZZw��F�ʮM!O⽋�vea��	߆[��+wo�J����N�d�4�7\1j6U*��5B_�D�R�*�+k���A����h���O=�Q�e� �~�����"9� ��ё����+�Ƕ��w"mp2�E�����C�拋�x O��~o�{�`鈼�[.	��U!ېu�Ap��宣��Kb��>v
� {��'����ȅ%�zhI2��� $�sO�c	��G��i�	@]�0��O��r����4К�q7�����Y�r��m��n��.���[�q����wB~�E�X5_��/ѭ��$��4�~Bv�O��q9��9h�r��r+B��Q��(m�P��T������$h��9��U���$N�Jȍ��L�ف�
J�#������i����� >��n9��_�����'Rh[&Uυ�� ��
�)�~?���>٭os�E$�
��%.����� ?�]rÂ�}���S��b\ eE�����dm�g�U .s���7R��0ϸ��_�d�<X�ݭ�q�"(ho�TP�B,^����Y�4�&vi�������zb����8!�W��Q �yZX��2F�6�&Z� ��[��mN4eMEn�s�gk��+>k� �X�E .��'zI %*�&�v�Ѹ��x[�ͅ�|���QrV��hf�}��Wh��_e�`F��y�2NO뚎�oD�?��tV���vd�)�EL��Q��ZX$�D�M���Ђ�~��ܶ�[����F�������x�}�)�2Wе�2[�݊j/z����w;�Ѐ��{�4�e��x H~�ƹ�l.b�A�G�|�H>�KMu��2���vC��t����!�5�U�e�����p�O0oX[',��R�K�i&7����|������4v��_%� �9Z�����f���lUW��n'���jrJ����\u�S܌�1!=���@ �v�r��^>�7��/ 0�Em�/`l���?��z[v�<�b~pC�HI1�����f�����b�GO�X���F�����@Fu��!�X���ϲʹ�ci[����3�Qnĺ����F�7���O`�{taH�{�Iᱳ�G�!'Ƨv�����3�D�$�@�w͍p<M'A�����` W��e�jm~o^��K�I8���Cm,�����۪�ӪC�)o�[8��\q5��3�յ�%���}��s)Do�K@�Rj�߻�un�zu1 �Iۻ����;^7�XkV'�<����
������̋:���]�AUR�'9v����|�I�l>�=�`q̯l췖�Rt�n,�,�,��EP3V���'2�am���+�I��C��1���l0�ۗg�N��[�,!�;�Kw��$WmtA��\��^��2c�<b�D ;������濦nb�6Ƣ��g�wkU������{6G�8}��o�7�[gÎ��k��
�;Ay  ���kf��A/���g�Ӯs0np��^���� �v��5?R)���X��߆����&{�����0r5��5�Uv[YC;��9�������(]A�d-Uɶ���`�A�7�9�L�
�+Է=Bl"�G_�N�~�&��u�/�I���w��s/���׆F�?�h	�M�+���H��W/V���vH�$�9�I�Z52aǡ#mE`�F����
���D���8����F�<O`l�Xs|AOK��Y�^rh��^�\�Y|��N�KR��V��Ic���:���wE�D�t�-��\��A¸_�)v�Ӝ�j*�����/߾��	�ͻ�@���6rlH|�2�PCE��*�������F�]�JI�6��Cǩ��$�of��ES΢,�����]�X�m���΢G�(,Mi�-e�4�}O�ÙN-��������u�� 1���F�`e�4�¬�5.�i�)�ߕ�&��3ـ���`��d�v�V"1['Q��FY�G�;)T��?]�M�Kf�Y>Jn�zp�*w���~�(��)� h���  �R�:���gAs�]Ȏ�����m:t��P����8�}��ۏ�Rgk^�c�_�)_�����L�j7!�/���3�=<�m�k���;q+y��&��|�EeT�U�c<3�o�����8�T��Ƞ��������n+�`ª�x2�,��+%�G�