XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���8��ݚ9�9�`����Fx e�l��H��j����oz�yR4��p ��(��@^�t:pv�;i�*��/��ބR��;�,�zt�~A4.3-Dn�BH����v�[����4�ظ#"\BC�斧 d(]M��eD�MNX4�WB��>V�Q��ղ��:�F	3�I!�#�`��:c_)Ꞽ��u w����.��P]Ϸwb�ywȣ#n3:�->���~o���y*r�Yö �|˛y�z�c�C��8i,I~u64[ĉ�y��\�����>����N���)����&��˾/�n��k�l�xr���uߌ�5FFq��6�f�a����I`òàȼ����~#.��'͛�/��:8�'�)o�����c@W�y;uQP�ގ�k?f>-�Ȓp4�U�H�E����$��F��'xp+{S0g�`y34P�ߚ5����ޞҍo��ӏ�/��v���}�����"��&���� "`r��]�nj�ͫ����vB�)$*��Rs�@U� ��:�^7�����Ӵ�u�U���������J�,ը�������^9�x*��8�� jTQ��3��"�?y���$:�y�|�������O�t( ���6@�E�.}]�́֩\�yxQѿ1k�xb��ѺP�x�X<i�I�C��j��U����p�2<���vL���9	0*��`͌m�w�����R�`i;��-ǁ�N�>��ʹD�$�c?��"��QvJ"9bD�j�=tYJ!gL��۵�[��&XlxVHYEB    fa00    28c0Tã*զ�=?�_�
�ߌ���5�L�� ���Y�ʍ�m����Z��֦���
	Tf:&)A�>&��W!�$�L.�QQmם�
X�N}3!?���޿�A�Ҏ�D�ϕ���z>�A�*&���&O�.���Q�����x�����Wd�Ň1t���qү͒�<ӄ��:����l)	�q�n�P�Ƶ�9AU�NRT�U ��JP%�c{��K9Ws��{�OH�!ϓh������ߤd�pC[�b�)'}���[�r�Tԥ���|~\�a��1��	��JzD���,�"��ne�b�^�_�&�\ZU�7�t��l0�ӷ,c�N���l�{�c��u�ʊ}�x#o�e� z��N��8I��y��}�,�U�Q�a��pj_��ݚ�K�> �P��	ҏ��/5�ň��g՜�$����"՜9��&2|a�ԅY8 ��N�CE���Ҕ�-b�Y�
tz;�h�w�Jzwؾl���ͣUa�R����2Z�c�tッ$ ���2��}c�_�j���ܦ��y ������Ѐ��mnN �ٸ�c����O{�lߡ����pR�Pv��Z��	E�'v7���2
��ԯ��eˡf��:�B �!�	Td�p��sS{/��h�B��p��C ��>�K�m ��4;�g}���| ����ֺ��u�h��1/�E���#��,3�85���#4!��;����8��]�)�p\�^,��D:�{4���{[��3Vtr]j4�&�a]�}�n&v����&E�*\|��Ev3%>�bF؊��%��Ď�ە�$�:%1]a��]J�HK;g.�,=仔��bS{�ǺB� uf$� 'ˈ�d��P���	��ǜm,B���Ǝ� w��ۤ@LkY1�H�b��[NO\yI��Й}d��&��U@ht� '��X��QA�)"WV��|����1[�U�Ьd$p�ޫ@-��EG�+ 3|�ؔtvkEg��0i�����tp����f�%
�l���=+^b�1��TL��G�n��"�犈��9^~,�J\�`�U�%,�Ta�9Z��JX)b��Ո�j#Na{�_�p�V��F�I��Oy�#f�8�w�,�~��t��70I�p?�d��O;�u�LF����99!b8Й��f"=���-��ʌO[xzG�F�SF�M=~L��<���4_�F��ć�Ҫ�z,f��| �M���J�U�o6X˱��j����R�d]~MˢA��0��۞�u�M%���$�)��.R)-4h�iO�]Ŭ�{9�(n����0}�{JjS~D��@���1�U��m�ص4����bu�������[�B�B啗��r9�4u�MF`F�@'Tg�cMΥ�r�66�����o�+_����J�fh���"t�x�I�K�G��D5��,�E�7Z�� 7ۧ�k�'FI��,��a��S��rׇ^���#�5�X��Y���y�Z�9u�^���Lj۰ƕ�t�Q��t{Tۗ�5����^����	�E��c�I�  ������h��8����"|FVF}/���\�Z}�G�y�(43V��]��Sw�b��V6 ���7
C�f�5) ��8�U �(g˭نb����c�l�审[�VqX��ՠnD����Q@�=i���Y���m46��O�ٕ{�f�J��C��1dk�� ��q�>9��47lѧcu�����z��	li��$�`�Zs%V>�6�z��uI���=�(������š)���BQL��]���Pl��MK���s,p02�ӊ8(�oo�>����:w��u���Y��.�j3��p#k(BS�>3tD4�}���NQ[���Ԡ��|�;��b�)�۲�Q�g�h�v���s�ס��V-FKM�����U� 0�L�c���L���"q�c�w~䱬����:2xu����1�"�R���
��v,�Q���:7r%������hP)z�r��$��c61�K�RI /��6�ek�ށ��e�W�'��tT�V��@n�ɾ>�n`ќ�nKD聯I��H��t:<�ߖ���v�@Q��H�v�7F�j�[�#̊t״Z��Գ�>q�{ /��S�� �X�KoꗋJ@!���Yw[=pŸC��]68�@��ZÜ���H��ةo�8v�B���@��P�ni��f�m�k���F��9��~�/�7�[C�邺��c� ��S�1���?;�3LG�CB��n`�Gla~���G��h��;ݞ��OB�Um����&]BМ�< %1�x��d�����Q�Į�T��zc��Ԗ0�V$��@�2r�Z�&܍p=5,}B����=о���h>���F� 1��l6��qD���w��bLԧ�Q�Aa�6�� <dN�y��OBz���wX��ڨ�DU��Se4�c)��"P�M�m`9D��JZ*=�	�-WK��v(v~Y5d%u��*8v��D�2\5Sb�U'�`��!WA����%�q��S�'��S��Z��2���L��v�:��2��+m�eF���2�A}�(���5W<�p&��؄[��/.�����q����.(����6/�O���H����/����>� �%�h�]9+�1K�ʺ�u�ϡk�������]��-S��b7t����^��"�y�� �~�p�Lǿ�����E�C��'�����?���_��3��~���Od�yqq��r���妒���G,S�":,	رϺ��!�9S�/Bs�/j���1�?�d~����4�7Y�)|�}U4kB��Q1f�[�b�/b�f�Jr��9�0�:�A��8N�nԂ���K6�Z�E�cHY=/����VvQ�"�X BA�l=J�b�-�ɂk�vX�DA5���t
�%�O�{x��Cu�U7�]�ԡ�3��-��t��Wǈ~���8�tFOn��ǐ���u���b�úH1,;.Q��f(W��e�.���z������c��}6b��)J���I%�})�ù���p�h(��e؏�s�%��!J~�cvp�A�8u��s��p�g6p����.��4�������(�Ŭ85P��>�#J�_Uݔ�e�Q�Ve�6��)�c��[�u	��P�X�j�4�zPj�:� �oі�	d7�v������(Op�t�:˻��1�c�G�NL���9T���9��h�0v~~8����'+�iƚ�fH(�X�eai�HUV�C���jK�j��~`n��	 ��;=���ݣO436��+M��@���d�3YAC:�!+:�R�qM:>\M����5Șc�ذn�wn�;ٖ�R��y|��,��9w��ӥ%��X"9���z�9�[=������V��uC�-v��V0$U/T��'�
٦���h�_����V�kL�EK��z-[u;��gMjul�Ze�J�造hcs��\��B�^���9,�c��'֐������?�=$_��g�TCz.2�?�9����ux��~�\�[�_��v^;pdԽ,��s�I#�3��0���"gߩ����p9��
�>H�	��0�V�5;r����)U`�C~���A�̴�Ј�؏��E�#N���Ѿ|#�@��O��1�H�5�'�3VW!G'� �b�L��Ѫ���/�t�/ �m��~9#3�Bq�-B6��lm�2�����*��[;:�-��ۧ3�W���yII��+>��A0�n�1�֟�ͬNMVb���_H�	�{���p�9k�v��ķ꺍�wb�Ӎ2��i��P�ӈ	�-�&|��O��&-N�% ���h����g6����R�T*4ߜ���=oe	�� ��F��؛��C�I�{����1 ]2�e���p��)�݆����[�.����_���f�O����s�����ne9,�~0��Cc/�JF���8¨���}�}��ó&�P����%�-!n�~�,��8�����4	����aO�����j��� ���6s�u�&�y�g2�TZ�W�v��7ڲ&1��Zf&�a�������ס���j%gĠRu8>1,��RCѧ�HV����&��`�&�����73�@/�φ�h�w�������)��d���?�Sᣝ�(gJ4L�������+Gu���VlۮMm.����)���g�����Ǔ���*��Ea&X��2e
�9�ۀ��o�k��~��
W���%����B�r�z��5��7ѺSR�.��'�;=�9�O��Uċ0�'��S7���g��W�p�l� �0�XWL�8T~����v�P읹���Pl���s�/}������o[-�!�?$���z|��`>���o�H��}WyV�5a��9���"&'��9������!Ԏ^�N���PJų$ۜz�O��_,#���Tk\x���4,���Kl1H��GH���=���LXxi��O�����ɸq��8����\㑻(p|�u��h����Ry���J$��:��>`�[�$jJ�?�õW0.l�)�J��C���婺&6H�~.K|�[�C��UV}�p�����s�[�
B|iy���� P)�9��ɬ(vU�@]����HΜ
��a!�E_"��|4���j ����?J�ʏ�T�f�|G���kW�Y��F��4E�P$��w��'��*����:��׷:����%�{�5��`&�k=�M��3�ڪE{M-S{�;��U��`'�V_���K��G�d���u%�ç��"�z*�J�9b���vY��Sle����3yG�V�&L{�tD�2t�zJ�4$-j����QLr!�8D�[�d��w5eQ��W���/���;h��4Non��s�&���L�jbx1�!���70)���<��i$��C�|A�	���c)��p��,�N+4�)��_�5��0`�l��c�(5fl9�ٟΦ��R؛S�"+��3:mZH@ڌ;&��4@DtO���_�+�7�-��D
 �6C�g�V༾��>ۜ�U}�k�	9O/򅌉g�&��d �%�%¤�9L{"��R�
�G�1�#z����lkU�-R�pkq2��`�ˌK'_�č@v��(3\�Lc�vH�p�����	����b�uP|�v�@)s����m���~���y9�Q�=6X��*�T�ጔ�;�u��P.����K�f�®qk����=�.-�l<p�j�{�e�Mcӡv�`Y񹕉gG�����ؾ|�:@�.�8?5���p�I�r�W[�ݐ�d�e�/�HA*�U=�`�����>ۥe����|-��]XY}�!�����B���ɨ�78�����و�Oc��]�z��q#vlI�K���� `Wt1�񙙒�4�cP|"%�fi�$���M.O�ހ�������
t5 ���jˮ��* _hr���G��WD��ܭ���P7������a�V���}uI�-�Ε�Rh;KQ3_��a	����#����P$[Gx�&$��\|����U?Dnv�d���~�M�A���Y�7fb�F����G\�5�Ǝ���{�9TUc��zP���)%1�����{��j�ɦ͵��DA�/n���O&c���K�ίǫ[����<�m꜉=���c`��]rZkQ�� ր�o�w�"ƊB�L������H�!b�-\����&�i�/SR�Н޹,A��P����j1�{��=n#Mػ����z7Bđ���D(���� ?d_��Q���=�mx������o�����w�%lͦ5FT5�Fи����U�,��O2��I�O#$\��b��iY�����"�����ZO�T,��3)����%�x�&e�H��Ċɀ����9`l�z�������h��&ybA��.mw� �zw�㿼��|n8Y�(�ASJAvMb���{�=��
f���̱��m�F�Zu�-[|��W:�<���l�ӆ}���γMt<W,��Q�Z6;0�s,c��x��9�P���H��6��k�$ڢk�ǕFM��ū�w�d��<�#���U��5���y�p���*S(,����R��|%Ku��
�� ��U����F���9�W�j�[��X�=*6�G$�W���l���v��J�^�> [��D������vF_��ea�OhS.v	���B)<�#	C)����$�nY��N���Dި��Er^Hh0<�L�@�4<�O�W��ѵ���JB�⤜�­�S�7"�`v��W����;8�3u[�Q��#T�Y�8��_]H��nH�.y���?�Bl��2����Ӑ`���(Rන2=yŎ�yq��U!���Cۢ��'v]R�����.Ĺ�Ý=,��1��N�%`ϱ�z�`�>�i��[ ���t%�.�)���9��g���i��ĕ�&��������D�O�cA�Z�hS^\����'JZ����zS%�
���&��46D�梋������Ami,���|h�B��la�Ѳi���7TUA�&��I��|�)���=0��!h�+)&+�����ؖ��a�c�^�0 "0���T�t@�~'|�J�����hLt����:ѱmdb��Ǔ7�F}�n�M�B� ���c��SX\�,&^'���T4m��9p���Nu�@�9�_��~��Z��,	�}���
d�
�~^��@f+=ǁ���߯r�a��s�c�h=�AH5���Чиn���Ɲk`�����z���O=I��.����$�tJ#�j�����d�Q�-O/g��'o�� 3$C�7��ثx���}L�͡��G�q�q�n���l�4XI��6 �~�۩W�E$Y۔\"�L[���k1� _`, �^F|>�;ۆ��٣n4]���m�$ok���u>Q��P�(&ķBc,ۛM\ƾ飲v��~{�mU��}���Y!l�H�b�c~�%�yNϳ�Uru$f��%)�y������)O@�j��t��je��	1K����j�����|��߸�E��_b���o︾�* CXD͊�Q{����W�It ���Vt�u����rt0���a�5�����|�ȞB��O3\9�4�&7Ď ��a�@܅]{��)�4�� �4-�I��@��7��Ù[��ꍘ���8g��z߇re!.��ԇ�mʼ�[�G�'��pc��C��VN���N r�5�*%"��lu�˞3�>�XB�6oG��ugœ�<��u��¯^`~NC�o�X�R��v�x9��`#�!#O�:UB���0s-�$�ph����F���N�)V
o����"�?/H���F�O����~"�z.)d���b�A�%����������	�������ade���+�9ւ���JXԌ���v���ͭH�̤��f�+L{|�4\�k�v-�_�)\����`5�}sW��0���.��9�w�!6�}�"/�^8J�@���9�m4X���7	���mƨ60��\��!of��:49�\�M����J���ա	ヂ��G��I"�=���G�y,�2r{˓W�X�04ϮB괕���/@�.��N}�{[��� ���å�u?��%~��c�Y�iV��e�{%8x0��a�,������PiT���Ж�}�33�e�esЁ�T)��A0��A=�*�P �١Ұ(.Z+��H���@��a�Pe�-�FGdR��BQ���a�֟;{0A��⹲4/��%�~:u371�MLg7`ů(Xf�����Rru���~��V�ix��X����%N�Xag;��'��"�x��1�O5��I��������L'y��j��M�눬Į�M��_U�S�ę�]ާ���@�7�eV�m *kafX�k����
>$��¾V�� W��響ly��TtK�� ��9�!@W�d�l�<�>�t��ic�f�[�d�eRߣYR��3�d�e��U{�8-���S��}�F1^�rA�; $�U�T>����]򑷻A�K�p(��K�h6��ʼ�r�"e�6�:�E���#.��(����d�]�bK'�k��YAT�*)<,0o�`��회�؉?�vw��*!�����ֺL���/��d�}����T�������*��zmKW��O}����؁6ȫh �.�5�	l���n(w8�h�5Zh���?.ӡ�G��A��}4�|��l�E�e�p'��M.L�m�p7��d?�|I5�x|O�fX�z�?�ج%�_�t}e�T���Y��� T���)FR��P��ac������U���sG�q���í&���9��<�p����O� �8���[�7s��Ƙ�$sz�Ҳ���P�g�2c��n
���-Ӣ.��bv������u<"�%=8�o��`=����RΑ���F[rRl�T��� 3���"��3 ��M
u�N�x�`�;t�N?�7�|��O�d��d��:���F���^`�l�n+j��@ǪK���'gR�
 ��s�F�vm�X\��Ϥ0Y�LZ�l��e���|��{If�����[�Cw�1����f��u�p@0��Z����C��1�p��SYU�A�6��ۂ��O�(>q�0�M��smή��Y:p��Ҕ#��I]X�mx�F��A{��Q�Ӿ
�\n�����
'6W��������<�T���)���V���ӹ ��ԉ���6n_t�Wڳ(��mlO��$��phнC�cʅjQ�9�v%:��ս���2�5J���=����/W��}�[�ɨ������M�̵�遪������di�^ b��	�Į���=i� b>�&h����)ۆk�\�ؕjU:9/9Wm�k�#�	�A��U�茙�Y�$$�џ��N`�Z��t������lYF����y/|"�H��p�df�ej�c�u�r�S�v�`��)��z��EL�[�q/9V#�/��.��h\!dB�����j[������
4�#���y|_.�/�Sxm�ƀ��3�Wa�S�P���UD&w���'�ϵ�k%bY���17�Ն2��h����\�S�eʚ`e\-��c<�Ů�t�.DMø%�N�p(�C6<̡/���ҽjy�x�*��I�����I�'�|8���A��S:WԞմ�S��;�!8��L:����dg�OL�*�A��\6�
^|�4uQ{�͠�%*,E�K, �kŮ��7f�ƍ�����_d3
Z1y>r+� -�����m�;���㟿YϞ��8?9%F� �L�ܙm�Γ��5�>��j<7�cT��Sh�Z#����q�ۧ ���n���M@{�s+v,}����p|�A�"�#�it?�=���V)��Lx�n[�Ο��6׹��|=HV�ap��MXWPj��.}�C@��1{{��LԽ&��2��)������f�=nTu����?0���qF� =��%c*�?�yю�x%]_�?{�,g�D�b���9�^@�	�fT�e3�ϊ<*^Ѽ�5D�� ����<ǫh}�4���,��y���e�(4���' �QϞ]�	�h��L˃��s�z��z��w�-\�R����I��8T���r�� ֌ۢ��	�L���y������2�{nÃ�3t/o3T�%�S������7s�;{'��~VF���%^�֨V�{I�����x���lvyߙ%^)�+����0u�k�u�U�k�)W8���f���� �꡿#�x(�zd������� �V�v�+b%��<Aj�fݺh,�l:m�{"����w<�1P�z_! �>G�l$p�a�lkFf��I��{PLE}��6�m���5��˳Oe���%�$�|�o�㠏�Z�s.�����_�0|="/:ZRq�����$�<��4���0�W7�Y���4��+����*�6�]*����#�W@���#�4���ф]�n�k�y��ܯ���J6�\�*탫�<<����=��Pݥ0���i��u��UEP�p�߷K�j������#M��`��|>�97���wR_���);F�,���Ҟݎ�|��:��CF5��@����H�}Q��/x=�˩�x�������	��1P��*�T�����'��9��`���ɔ��ܒ���,ɏ�ܧ�������u�g�Xh������S����
PM[�z�՜��~[�18"���z���K���M�E���	�D��yi���<c�)��_0M�S P�]�����1P>��$��8�6�LA��)��ejAl�4Z7�~^�/Gn[�����'4�9x����)�ʧ�qkD����)L6�<}7��7�l��uXlxVHYEB     896     280#)��GmJ(|�ܛ�v�����q�)�P�D�>A��T�MY���G����!CR����k�
�\PϺ�A_�م3�wl�_>�E�ؔ�@i
�e9w\Hp�<)�O`��_�+�R;�r�T��h0%� ����&o��]����Np� ޜQ�$�?�k��u���}<X�q6��)���w�2���!�'!=��E޲^}8��W�_M#l��$�E���"g������?LMH�	j�h�r3�#�8[¾��^�+֕:�n6��m�V�����]�y;���I7Q��V�n����c�TAD�7ϥ��ʀ���e$Tx~-���b� ��1�
q�+Ll��^l<k(�ɓɘ���B�X��*99.�(7���Sò�m{�6m�f�d�x"���:�8@m�&o?/+#�S=z���G^�4�R���h
��"���$�t+�jiʕ��A�7�*��rɦcT�����j��v��H ��퐶���Rr2��׭<�2a�rLK���g�b�D��L:���4P��n�;�Sx �~1x��	QЁxuK��Q��� 4����TY�4��a;o��äq>��}�üZ��Fj撉N��wN
u������Iye"�?U0��L-c`��3_;�����7�l��ڗ �Uu�