XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���!Cs���� ��/y�+q��)g�SpB���k�ݎ)����%��F%E+0d���s߶o�WR0�;�@
G i^�w�OJN�~0��U�ʋS펕��i8;A��r:�P���)O&a׬C�\�T���&�@�8��e��k�!vؒ��Qj!�9�#��`k~pk�mt��ν(���5NJ��"!t9�'���ҏ��m ח䧾�}�"K��L���� �xEJ$q�f�D+%�%c�P��y;�[��52�w72�k9��O��g�sd�[�TX*���]u�F�q����'�!nK0PQd�D�R����B~����̊Q	��?���1I�a2�1�Hթ�K�K�������9-@6�&1!}pY�b���Ն���ndcr��
ay����`ި[�D@Em�`���h�.���OT���P�v�Z��գ�/E$׽����Mr��bE�s��Vn�w��'�}��M�I���[�,Rh]I�,7v`��
"��/�Ѹ�G�J8�깞!��=�:��ld$� 5!4���K{������a`��h�#����Ԡ��E�c1��rr���l���K�?7"V���̈́�����s�jH�?(.����[�jP#�0�R��p9�Єޯm�i���؇���Gж���y��C'�TFv ��2�֍��M9G�'@��e��m@��[b=T�	u��B��M,�& ��k}h$2LB�����#�+IǮ���A�6A�;Ň��F�B��XlxVHYEB    fa00    2520�,kq�Nd�\���葍���v��@�OC���D�N�U&¢$��B�v����H���D�C��now7�*�� �xS"]�.1�c*6��oa���C ��[�H����I��S��}�~�,�T�s/uf�l��<4޽.�_k$�Hb�4� �%I��4�ɬ�p�gC�,D�����\ni�$�@`�r�t�l]�||ƮC�H�t�mʓOF�{���׍vP˹���J�t��iq�s�	yi�k�P��Q��Q���=�7ݯ�j>���ͭ�6`j��^�����D]Ո,ō���ډ)9���4�{���y�m�E:!;n�;�$1�#@��o����SF��9��܊3���U����J�,��?m�-D�J��&��m�^��-m+�h�Z��%�$��66v;׈�
���?���y�Ą ���o(�0	��o�o�X�e�Ĉ��\^�V�@)���q��wM�),OP��W���雋�a�D�bZ3}3ޭ<Ҙ�
�+W3�\�N�;w�DxE^A�n�I���
��S��ge5ؙ�-�6 �h��p�Խ�lyr2�m��i��ђb�G�H��J�����kЏ�$�r!�N�~��Z�;D��w�ϝO�]z��۫�a�Κ�'���J�<���N�9�u1!7�@T�y�V\�*���``~���iO�c���>m�
�/�ҘMb��!Þ�'r)�,fLƿ��"��	5�3�����=E��g_�����w���&���������:����#��L�\?8���֤ϫ�\,bX��(�B��p#�yj�߾�H��.�B�p͍>>i}��6cĝG��-�KۛVJeA�MuY=;d����kef���ƻ�����8�T�mo���5W�,'̘B3>r)�q��3'mt����}�7R�Y\�Vt�r@c'�5F+sz��)�U{�sf\֖���=�B��^8e� G�h�Z_|'"p�Ƙ}wp ��3�U��Q�4f���IW;��SE��m��b��#�Sŏ��-Z0B�u��0��U�Y� Ǯs,��H0 ���4��`�:�<w�4bB LG�[C<�z��Z��ͱ��=EE�̭�n`%iF�Y�'`|]\��6��S�JBj��� ���P��C���/�U��4Nի�7�^�-��!�r���\��-١V��:��G0���+�oQ��/:�H��,)�$�I7bT1�3�fC!�� �u7�c�+�l'o��Z�x�}UM���-�����Nf�,�.X�x��B���y�/\��Zt�`M��<:�k�i��v{����h����M���ȣU�1�?���w4�7��LC^!���ķ��F"��9��т��kP֢�����w�6M2큔G:5Ě/��Nxv#�[����`����Ȝ{: 	��T�b6�&�QiEE��e9�v�-��ϾK
\��=����;�k}�Ib�M.s���zTu�n���Rv��
���K[�;�6gPn��E�$'68,K"���uQZ�����R�ר~��H���~I���b���`�N�?F<���E��_%i��]!MG�ʝ٘	���I	���)��/s�쳌�����9�OĔ�f����>s����Ǵ���
ܳ��z����F�FAv���I��Ixў��v#S�`_C��n.��}2Rz�$�q=�A+�c�	��.�]�ϓ	n˘��=�rѸ�q)��ɣ;�9�|z�0�`�r��'[qm��F���$+]G,�����%��zKBY�4�K�����ZS����(u��K�j�up,9��� t���/D;^�gc�6���k�"���m=,ppe��g`	&�e�.>.��:�� $�@D]<_߲��ې��ѹ4�mN���Q(*���z�q
ӳ�$�WF��'������ ���r7�ܣ�iʼ�I�E��B�`4M��=����i^����[����!��A���DDWpR�'L���(��Ad=�Pci\E-��~R���v0=DZ��m��R�&��N�O郾ʁ��W��H�2B��:�۟�uY�\5����E�Y$� �(�B�8��-T���F��|FCR� �o�|R�$k����,ȓ�{�k�9{\eYl�	>N�|���\Y/f�_E�P&��\qgPU�������1��a�ӻS�K׸UV����E��=Sg#���ޒdWv/2Q�3�xٕ�i����HK�A}2��ާ���T2��##:���a/Yۼ%��4�1|/��!��'�Ru�F]�[�3�@f��NSj�� �G4�Z��"eUӯOA:���JE���v�8j��Lߑ���)�*�M�,�7Ǡ���7�����7|"9�TPӂ�����4<܁����k V ���ɭ�n~k �6�KJ,��@�����)�������(gUw<Fc{�S�8��`�����F��~�Xrj���o�Ɋ��2EQ��2o2 �5�>w�Q��>��H��������j6���IhZ���G�̤��Ky�Sj$���3R����zv(QCs�zʇ�3}��Sb���wi�$����3�X� 1��D�wGe�a�w܋�;Pѓ)���/�:"�1�3��&���>�X��uNJb�.l�M�|!������޶���8z�'�9�*<^��T�\}(�.KW ��ٶ�h��w��P��T\�ZU�/J$66����<�����ӝ,�p�أ%��i*S#Nmr�N8z4Sc�y� �Λ�9X�����{)~/��\ (��261�'�8O���TSI%���8m`Ȭb`��z�z�c>x��b���A\W�8�I��=~Ÿ?1�FI]f��׹��\���#�Bm	�L����,c8���%%�����{2�p�����٘0���p�\�w�l��)��̺�H��gci�E[������/��j�$��/�!���g'�^�U���~�~��*��抰S$=�4��H�[���Cı�1v��Oǋ�j�ݎ�ck�%*��uYL�7��M�
dC=�-؎V�ȡ!y�t;�ӄYo%�)2Z�6��CC��
�@�H�L�W���eBa����/8���s�\m,�ЉX��a�C�%+~6�7����`���$t)�}l_cb�]��<^��`��aY��D�%q�����*$�~Z�C�a<X�W����	0Y�z�w~݇��8M��P�M�x��̄:P��HK�Uz-~����-����&?f������x)��~<�-�?�|�+��>m��)^ƒӗ��떘�tr�8Mh¾<�
-s�J�m��o�Y�$�J��lG�@�$�s��;��2UI��Z���mx�>��+c.�al�3�\�UCO�-�� "��&��I���U2.2Nˣ��1Ћ}�N���,��4�>|K�����mf���@����$�wtP���\�.Qڷ6�B"�y�����d澒p��O���9�fP{z�S��'�uM}ܪZ�ݷE9ݘ璦8!Ւ�5h!.bH,�.��B?�g���|_W:x�b�D��;{����q��誛�$O ��+�(
'�G�p���F*�k7�\�ى��flV�F%��q���/�����J|�FGH # �x�Em@ES<��b�N����:�L�=|G �<?���d"���ER6�8JxlɖD��2�N̝���#��n@�$��Q�('_���o�e�oF��	i�_��k��]��'�2��ŹA������8s����>K'�g�Ml�<�,�s5�:��·4`�N�$�D|����:P�����摗6(���|�~O�c8�j-���piu�y"����ݖ|��gbټ��l�ՄҮ�V��Xo b������)�7c��s��s��	(����>�^d ���!hW�w�&�;��&���)�}M��p��D
3���]��|Tz��"�d[�7h̆`8�/��+�o~�M
�M	� ��֗�LJze�Ѿ���.�����@zF����������+�l��W��@��4��5�>��B�xo����`-��S|LK�<7z��=�7D��P�u���`d�>)L��ک�2�8�y�.���#$2�2�~�ӣ�S��R�W�,����E/ŲŊbv=-���}��i]SE`Ώg�-z5*{]ÁJf��mH���t~J���W?DL��yTK:��f��}t]��E`���*����b���E�A8�"��]���x-$$�1r��':5��T��O&��p/���o���]�D�8|Q%�Lb���4��p! ���@����2W"9��^Mh�ڦvT��`n�e'a"��q�Q-k��gb'!v&1�0�K][��	�kUV�>����-:9d/�j1hѳ�*�ur�ʇ`]�֛�]B��(���\>Qg��% ��а����6�p�k.�PG�>�w1Ὑ^�h�DGW[�|�L�4��R�	޴�
�-��I/��6���sj�yiw�rF5�6�*�82k���14��;�;7�:�An��'���<m�ǆ?�텥2�.�s;2���=��d�����w��:�дy�) �T��`)�d�@b����|//�pmی�����^�D�y��"�Lf��Dz��Į�Ew.�%���w�L��WZK(�UR��x��C�tO��&֋������3�3wMDD4q5ӖIk���j���99����D����-��h��nc�M�a�(�3��jp�J�<�M]/R�ޓ��������qJ;��~jӥq�2��5.م�+�����A�6F~;F���j��>1�1vzTs鲉�
�46�+���y��	�@�wt*��%�����>�:�j�xឍ��c��6�eBf�]a�a����t,gP���X�2����Eo�_щ/���o:z����<~}�h��/��(e�L�h�8�4e�N�BY�"����d�ut�?^+_A�yL�O����0�vý�#��Ӝ%Y�b� �q��4Gd���B|���Ǔ;����(� 5}n:�uh�|���=K�"�U������cɨ\	�r� ���ͮ�p?�d3d���\��E =�X��H�1{ye���Y7�.���!�Sc�J�On�W��!����U�ҐK�8�-8)�A��s�����è��_��yy?�^��GX2���%\X{�\�w�d��`)�@H0d�=���=d��<��z�9�����A�<K�	�
1H��œ�"��J!k�ՈrO:��ݪ��xL��h#r�����K�,}�����"	�ϩh� ��Y���ڰ¶M��}7E��&���-qaq�5y��r���N��)S�-K� :�P��3E7"���ޭ����N��2���!KH�x��T{���~�/EV���T�I�	���"=K�+�q��?i�羊m>�DΤ���E����i ��(�=��1�zv6b!s�h�7_d�<sH� ����RY���	��� ���'e�V� 1�<l���3�������y�������/[Uz�<�ǃN�2;U�pb'���tX�Ot~ʝ�2�=�؎?D�"���D%0�[�S�;<m��L���!Ha��Us(�?QT�c���g���<�AV҅��<�0�������[4SpG��Hi�o7�J7�U��7L>����g����"�8���������C��K��}�,B�ܦ�-2�IFlB�1�G�����$����uY��U�ץh�����7�8Ȯ��x��S��e�	����We/��9b�|J)����ze��]m�ӻ�(���HhѥA����eC�nB�j����i+�U��(��G���[cf����I��7ı�?o>��템�a	� �܊	 1���a�6�t�؊"��Ã���$���҇|Z�V��0/1���UІ��MI�Ri�Bg(�?�p~����=�
�ڝ`ٰFX���2��NŘŖ	P���!�n��Sai��8��c��<aQэ���i�b~Ph��ϙ�隱�[H`YCO�K����0����M�D]�lD��f�c��`�i�2�����Ps�DH)kTx��Bu�|���#]
��14-�7�)-�H����?,,�����[�8��%��r?v!T��煍x�[I�D�����x��	���O~N"�!9�^�W��1�<N;[Ej6�Wt��U&8>�گ˵H�:�z/���j�fiBp��(�P_Y�OH����(�{��k�14���s\�3��Y����0�*�t�c�Zz6?+Ѽ�8!.�%����xIrA�l��:�����́�v��h�έ�#7���?W�ZF��f?��a�$ل�}hZ���^q���[c:GO)5�v+#c���{�'6N����Im���o�|w! )�{��Q	����f����y0\�W!�dqCq���h�i�y���%t��O���3�4�zr��!����e�J�P�e^{�IyE7OwI�A�F%j1@�n��T@EV��\�4a�Э�4��zh���G���Q����m��%��;8�$�����{s�\1-�	�sK��/�2W�����Dr���w���2���O���}�ڶ
��L0���Z�l�7����^���BS��a��s�`���_�������'8�P693��o�@�O�]:r#������Sk�r����ϡJd_��6B(�p����U1ۯ%���r�_�m��c�b��0��CQ՛>�K��x�,�d�d_�{��!{�_�"���E���c\Zi��xzz4y"�>O>ǳ z��p����v�������5Zw��TpP�����ԇS��j�]����j�a��5ĩ\ߊ�%<RgWy\��JqҎ��Y2Sy�=��#b^A�� IB�z.�k,H{�/�p��xi���=5��7s��h�����-\���jHj�&���ݭ�H�)t*�	�|�Y���SkqS��h����hT3�����?/�{�u�
��}�t������['Y�C�kwE*�^��RF��^�Y�р���:OQ21�{�%W����Fʓ�k��9��x.�u �=o����]'!#y`��އ,�[b#ͺ]�/I�(0�@���-K'��w��e����B�'�{r�mA��{�K�O�IѢ(ߩ	X�2���݆���[ZB=ꨞ� �k^�zmaܐ�O	�rm��&zY��~ļJ���7��
����s<�y�Y�
���ca����h�:N��>��M_&�TTu����&q���&�W��K�i/�����!S�3�7��(��ty���ַiۨ�}�
6,�T.,Z�&�~�w{�6�́X�V�D�C�Q�p�m<��|B�,>i_����F)���*��q��Z�4��� �����F:\P�u��^sx��C�_��Be[8����]-`j����S.�\��[w�h/OV	�񾐶ۿf�qU��[{{}ћz>���mb��3Q?T)Un�6?�,7��~u�X�X�F���Ω��y��?�β%��_G��ř�ܪ$D��>DG kJ�/4��s��C�-�Rq��T%����܌��uA��'���U%黝���݂#2A�U�*	��@2���* d�P�e\!�g�hR�z~i5#���]h8DR�p��՛�[�{�
`�Q2�	�w���5��ÆOo�%��q
�>'��\�2�F�*��ۥE��`��x��9
G��Rd�O��}k�b\lD�|̂]i0Q�6�=�I�,ɡp��m���AJn"vZ�`�$J�ԄT2;��&m�����fy֝`s � s� 0��l�5���	�h�����F��5��?��L�UK��t��C]O�x�,|!x𗘷��t^�!E��gδ �~ez
�>*���ԋ�V�͖��	�����͊_���Vm�zo-x�r�)ֶ�`��}�6���`�[�����z�%�2�.K`'��O�3�׎�'�_\��X��%�k`��e�ύij���9-~����cE�!V?�:ғ�O��Qs���~�*j�����$�Z��3Wu�'\k���n~�q�������
lAI����S�^��-�c|��m�=vo@^�x�t*��3�٪ ��mN�YG����N��%e�&�+��?�l���y�o\�څ�M�XD(��.0�c?�Y<��.��d��f�t�$�P��7�^�HV/���I-;���2�۶�����
��J�_��o���J�K�wѠ!�O-P7d�	����L{�*���:J�@h�������|���H��R��?�h	��a�'=�Cw���Y^M|)�YW��w���(�����^�G38�t��J%�, �6��zL�H�!����p\���s{�P0N������Ì$��^���Pk\vM�qR�����Ƈ�������Y���_l�m���#�u7��^�_�߈�kAo�So�s���ǋ����2�$q�yw���[��#����:"�Ǒ�b��+�D#]Ix:~"�<gb���Q״��nN�p�DU�� ����l�� ��'�����M��ͼ
+�e�iЫ��YטlW_��ǅ����3�#W;b��.��&S��!��辐t�է�K�!��D�ݞK��5���L�F����P�1�@fn�1�<�+�)�Q����0MYG%��μah�G��A�W�m��A{��gŧ��I�T���ߢ�Ă�� �;�v��.�}�D�!��ăp����#�#�7
��AL��ZM�Lh�g�w>���+��F����ר�n�̀��aÁ��¶�>p��gN��a��,���]ԑp�Єߠˍ���c j� p��ʦ�bq�񰓧X����k1��KD$�=G,�C�VQp�j�O��� �R�N�<�|�U�����`��t�������۠[,�������:���=�>�vgM?6ͣ�҉�Km��Ň@����b�����y��R� �\8-�6�ƈ&�Az�)���2� U�A
�p�\C�������C�{?�ˀ�EDOÈ�7̓�\c~Tⱃ�	�r�bQ]<2�W`Q����a�{DS�@?�G6������ 0�����q�Q��'����i�K	��{���T��S#_���3��؋�׉��5{�L1�<{�9수y��ڞ�P($��/���F��+51��1L��̚8b��b�Os΃snt��\ϙh�S,	4*8�j��n~��M�z""��u��,T�(J���Ɓf/pi|��X���!R~*���]b�Lޥ�WB7���
6V�(�Y�Q�Y���Z<5�V��T�
�B����Lo/�9�l��8'J�^���~^[�(�R��1�Y���utGN�'�.YN���yڍ21I}�0q�?T�Q>o�!��]�N҇l���s֕'V*��nt ���X1���b�40Wf>��XlxVHYEB    fa00    13e0����0�l0n7c�Jй�q�1��n�sa�k e��c�Rkg�]�7�C��Q�D���e�H�Cy���\H����~�Y�e��:�a�i-s6�)v?;�ی��ä$�� $M�D����y�L�,_��<%6�#�
v���y*J��H���A�9�iv�X��KsH���
�CT���4��V�+ˊ���\,�׌�I��d�\/�o}�f����aM�b�� 'O�`Q�Q-�k\!�����8P�ήK\�G�.��wry��	�L�}vT.��g'B�0E�e�+�ƹ�5��O�r�l\��o���ݙ��gK�J��&�;�6<��Y*�*x.�mk�{7'!4y��pȗw��Z�8f�C��(e�=L�P��JW�̎b��k�k,,��A� >L���(J�7Q�\�c�A�a���uZ���y�:��7�?U:����?�W��A�J����eo�	��������e~�N���X�='�<\�eY@#"C	�PA]�6�=(�) �ϱ�7e�$O�x�S���I�X�*��<o�e<���=����wu�Ny(�q����ɹ|��7��j�ڔ،�V;5Z�L��=p��|W9�bVb�.�ãA�R�O+��Xӗ�=䆔��#s�����7	,č�+�ϡ@ f��ZiOMc���}Ѐ"�X�^v{���������w�?�և��`�BW鍹2_2?YЧQ���F��Bo����&��xOM�Ԭ�?3���`���1.�n$�Ԭ���D�����W�'�m���^����N��99��9C�õo�B��֑�}@�3��,�ڋ��lƧ`���R �C���n�0�����=�ᘸ��rn�2@�
���qx�f����s����n�i�r.�����^z���^���FTCV(n����OEg"]��l�aъe[�aGfz�q������І�ŷ��E:3#vG���mtBq�%��,R(�+߬�D��A[dKV�������CF��{yY�4�_R{B��Pw ��M��9\~���O�W�_�_��SFZ�'n�)��p�/�&��[�+>�ZA��:.-��B�)���f��~Q�sp�����R�Mr����_ߡt����]JU;�;IG9(���"��)�=�uo�������It�����WSH�5 ������y_�y�W���M��an�
[I&�p�ʠl�4Oόw��n��р7	=8|�6��l5c5�%� �+V���<-�W1�3�r,UO6��f�H;��LY~L;��l4�+Wp��B/�@��c:r���lhL;���G����@t��XJ��$�0cBd��4`�*gD��2P���F5�@ ��R^�OR�ύ:,1�l(X��(X]���ֈ+�2�Xѝ9�����"߄O=�%$�r��᣼�Z\$�V��~Rrrc`�h;�y�Mat���ʃ:G������x^��"B��p"��R:���<`�.1ݼ��S���B�и�y��u�k�rl4�B7�f�FOZ�d�AjD҅8$$�M^_�b��n�l0��b��%�
W`5��H��-�����-��o�&������Hx�Ӟ�>��v����HB2�S|.=	��{��i���=X#g|I��7��S&�^�D��z�{�t��)z]
g��!�R7~�/ ��M�P1��b�����yⱋy�qd0�&h#��]+���6�X�!�6#]n �*�'���d)��]�"�TW�ms�5�{��y�K8�#F��W*Q���h8��S�d���x��@�S�۷���u��nvv�4��>o���T;t�i��/i��Ίf\Ģ��8�]����T�m�z�n����Z�M��B�f�x-��	�z��*�H����"��
B��$�� �%ig}QL�{�ql�Cˀșk�����;��48�[@�6����]g��.j�;�A�zM���v�v����n�A�����ԝcz'w@zmAX7n��d��{����%Py����n��cy�4��B1O1���7Z�+���_�U��'�.�}�c�{R0f~J�.kJ{�[S�H�@!iNښ |v�&�,�')'8�~��� �I�r�ڃ��.�E�JCk*\�o�B���	lT�W�Z���헞/Z*���E\[]��E��Vto0��l!��0J�Ɋ5_�֎���y�y��3�<E���^�����I���;��Y�������_�ZZ8��r�k.��_y:��HI�����5�B��~��-�Y�d����-\|���7�e]0���C�-�Q�U"� ?U���-�^ǯ���2IY�50�?\��j�J�t�M�O�p��ѧV|���N����=��Xn`�/;z��I��g�*�;\���?Ө�������&�3(�\Ks÷�u,���-6��"$�m�+k|P�<�?�p�T~~�Y�,;�'O��0�$�8e��|AT�ǽ�y�N��s]�V 9��%/��9~�	�w>��|�Έ�¦Q�v-���X�:�a��s����@��Q�a6c�E�D3��Ԋ�f ��}�ӴhBQ����:l���[�ό�EB_�)}�kk�T=�0�H�N!�{V��R��:��V��g���cẅh�����?��#k�g�c����'��3��Ǉ�M�2N�|qS���B�OI����%������Oa�Y=�"��a9I����$��^A<�� �x\�~RR�L�L@�[*ӿ
�C�6.�WP�{V��5����"2�Z-�u���I�`/_@�4�E�P"=A����I���������Z ^�"�8^׮�LE��;g��yP"�xjq�#\YHO���2��B�:]ԲT�lXL� �+����8|�'M)�%��T���KEy���/Sz�{4l�m�<c�� T+�>���a���y�H�d���^��W�f���R*b��6(�`H� � �$z)r-7L>�96*�j�5�ї���r�������o���;�6�C+#�֔�!*��e��?b�e���#�5̥�ͫ������$�w$9Y#e�J�Q�?_�;5f��]����D��x����O� >��N~7إ�C�b��GIܭ��.�n�jˏR�*5�4��l C
�XI���[��T�K[@�A�� ��H�����lSoS� ��EI��k2��t;��i���_wo�yl�n�B�{�Ɉ�S�) :R-��1��=����/����K�\� Ķ�8���vs]����YYE��[et���_}�>Tn �V�<�ñ-�욉�y@�]��ήѾJv�$e��o`bщ
������}��.�ĸ���ZQo�q؝�b�$�?��x�NVR���9��($.��*1�3�L�_	R�&m &��[Gj߆]]�f����6C\hq8�6��F *��!�2.�"�?1�΍��3�B�����Z]��]���Д�b*�.7��PS�u��1���+�x�&ϡ��,��U���(R�~��;��6*�z;��!��������2���	���t?�`#���]	������'��<b�Ź,n�J���Xa�[x[t��Gd�6k���X1��pS�1�KL�>]:�[�N4V���u��X̉b��!T��ǈFn1_��]��8��$������zN�v�[85~���X:l+d9� ��p�n���Vϑ� �Ϛ�/u���;͹	���Lf=��:�E�<1��V��oz�Wm2^���e�D �O"�_�4ͳ<��]0�o�π#\�0��\�O��;aV�[�e���)���5�L����Y;�C]��8����!���U,C�z`�vK�.��C�g�+ѡ����kڱ��ܯ�H��|��ӳ ���g�����#6�,'-5� ���W#�	k2�D2E�����9�_�{���Q�j�7�>#� �Ǖ���4IiP���U�������� ��=��h��ԙ�6/]WUۖ{��*�u�6�=�Ao�m�Kh�asj9W��O-�:Z� �Ze��
"��`�=�2��G�|t�"�z��,�қD�8�}�]ۥ�
"�~Q���(o�}l����ڦ3�cଁ8ನ��y�',�*�F�ٔ�պA-$'5�ŐZ1������,��	W��*�{�nP<���"��е�i�G���8k#����������6v��F%��-$�ۥ~�V'z���<���=���l�]�6�ϝ=�����o�@��D2����� �hTFb���ɺ����=|�
�\#��B&�S"�p�	6�l%�l֩�[X )��It.[�K���Ȉ�0��FO�]*�� 5gm�@R��=H]_�g��ӳ�xoԕ�h9��ݼ����}?���v��0�7;�>��C0蹩�QBX�Uv��]CI^�n]yZ�үj��M~��!Ř2$��tq��}��Յ��p�k);���̪�K����^��M3y�Z�hm	Lm*~�Np��/ߒ��(���J!�	���*�������Z��pȿ|U�v�$	��h��`�K>�ܷ)����(_l�Y�����L=��&{���ȯ@,ir+��_�������bt��B�8�@7A�-�`�껪9d#M �o�a�$�����1��>6�yPd� g��j�ʵ�1[=���
7�"J���U�M�)�b��y(�F(�*څ�.��=�=R �4�W饶�~��{`��o�"g�n��o���W�����>°=����,�����z�-h�:/Ȏ����x�a���v����Z/�o�[n�D7�妽5�<\^ә]��'�%�p��4���`<�'AT�υ���0�e�d@��B��� i=^����9��o}�zZ�R�@J��-Yկ۲��P�)�F�(p|�y�YG	�� q��9D�J�-�J1�3�V,���;�O����f�Li�H��}�X��n���].�U0���wl�5Ke���#�}��s��L&$�5d#�s}*=�|R���n���2��h\r� u�ȩN�A3����J�nժe��I�&��^�O�1n߯�_�(�<��XlxVHYEB    fa00    1780�qo׽����icX~.�������G����׾|�H2Lp:�%����yvg��V�Y����1�{�)�z��2i�����7e�]��6c�Ͼ��-���������5A�*��Cv�X�z�7lS�M�RzY_x�#���+��Q�Go@?�ꨇK�He)L`P�7��hJ޴���!���{r���Ϙ���e�T'�q<a���t���m�cB�f�`�!�;c,��'�)+�5�X�5B>����Q`2��+�����;�yH���˙�3���z���}���R��[�K�6Te��Ì�w��^��i�Ȭ.3>��X$�-#@�h'�o�dG����;a|l�h�T���L^�ֽ�Ĝ�6:b3%�6x������������0�`i����&C�ǿ	�$\M>��Ah��Ð�N�X(c:�U\	������FHXZg]�'����r��Q�Ǆ�J�XqNCȒ��|H��ND�3U\�H���H��e����sv���
so�Uube�f<��.���8c'NOq�NS[��ϼ�~�+�=6܎�JDTF<��<�o\��/I��&��0�:^x�Q��I#�$�}!֏�W�T�}��q��Ǭ�-[��.�&6�d�H��N�ۻ%���?�g{Eԍ-^��s�6 ��Ҧx�*�f�V(y�?�zggQ�[��t����*|��q
��0� !֌go����`u�C�w5,��W�ƛ�9HV$�2H�y�]�  T�86�9�Y�U���jXQL��X1@���)S���y8��R����>��)U�;3
�D[�ǆ�B\��<ٖJ�SM%��G��*Å��Kh>�J�i&�\���/~��5w���MB%�.��ܣRvuF
%螾(#��:�<�}�5��ƈ�ڨ�I�r��9T�3�����-�i�ᮯ��jd$M��J�������t��x�%�K�Quw�r�#ׅ���7q��	VڅyO�#��)�����O������p�N!%,�K@�P�����\���˩y�~/��7��F�PoC%e��ǦA��d��煕�@;�y�;�603'n��ξ�P��h�㢚��sb�7@���7,k��i|�D�����=��E��(��҉�L|?��z+���p7����r��Q�%ҖF�F�Ws��8��'L�����z�k��|���Y!}i�B���VJL�7��鮋~&8MS��rԦP�$��Ȏ����s*$��y��>������v T�G�r|p�^g�e5��c��[��al�֚�0��H�(�~5��ݳZ���]�@,5��	ϫ:&C�$�C�YGwq�	`�=�����R5�����TJV�#��e���[��,����7���+F������r��E&��
�Mw=���O��g}�n�h���ᶜ��V����;�蕸��e��7��}sC���+���XP�3�(��=s�Ҹ�$�{L���vP�|�1.@�Np.+[� �$��K��uU�����}�^�8Y\ٻ���o�<���a����V�	�!��X�ts��щ/濨��OBħA�&�jA��2]Vy��<Z�q���2�Cߣ`�]�s�kMA�u$�t@��_���-& ��&B,� �?iP��Ůn��z����O��x�nY=S��m���`����E��@���5�x!�#��y�E�8�&a<�����A7jӪ��by��G��RY�j)�7BK��e5�l\R��Xl>3H�5���ClH3v�ﯷ�4���:����H�4�k[8S������x�ĈE���1���r&Q����y�{O�B���f)�c���%4ٕ?��c3�t�u�	�4���_z�2����pΎ�3�,<e���DW'"��Q-�*N):�d�
�~���t�x��BUQ-����&1�Z��$�j���/����>&x`��_��T<�#땛O�R��d'b�F��o%-�Kd0���G��}��W��� ���C���;T"�	?h�35;�_��B��i�~���pU{+0k�}GS�7%�3]��N��d,��?`?yD�M�����C�Ε?��*���\�H�Ln2���E�J���*�i��o��1�N���%!��]��+tH���c �X���XJ�|�F���!�V u5��SH~%�(��}�-�*��Q�~�̽�d�sX�r�
:���A<��ם�/�?��7r��W�w}�_���_�sU{����B"�FKЯаJ�ꋦz�lv��dP��t��$ot�^3�)����8ςnj�ɤ��[j��7ߖ���KF8����du��n�/�ؾRJ���p	p�F�})�^�C���5I�?p>1B�j��������������s,=7�Ʒd5��U����q �[�W[GZ�:�� u��{w�c\X�C�[jEuX���C\�����-�₲��-���(�v�C�Yt�6�&�_+�Tr�`qMe�,i��8`ʮs8�i/˕ �#
]���M�!�p�xd���q�Ӣ^P�ؽ�IL�z���\�`��)�d�����qc���}j5 �d�H��jCf�	q��x�IQ��@�|�G�O�?��S�\�Ƶ3��NN�� u̹����c[��e'5Ȼ�ZĴ,��_����#��� m� ǵ�ƈ��%{�Mi���P?G�z�B�Q�H�����
��	��H��[�0��;�^�I� ̼W�8��0'��7�k�<�~@&*�>��X�S�oz��G�@n�	n�v�Am�ϓ'�h�Ýk�h λ�Q�O���>��kvP�z>�}�SS��Y��ڰ�C+P����Ҽ��k��H��{8mj2>< ]���=5l:v�=�Ҹ�G�О�rm�ȴj�f ��Z�S#:&��o̐w���>���<��// HW��k1$z�آB��\O�����E���2�"ج�9��{z�P���=DB���o��U��������9���� }��9�p>�^��ޑ���;FB%4)���2��7�ɢl��*��Uن;�]+}�M	)Z,sj���F�����*���dB݃�6� [����:�%��O�p��fV�bb|�?0�A=�9��J	4q�9�&��9#�ƶ����%�vq-7�-#��-9�R����2�,���4o��T�~tޏ��J��ǭ?�>gxS��vي>m܃����@\��^�K(䵥�&�kf��)7ӽ WNH�k.��`/e�)y2̫�*���)��5������i��mU}m%���Y�����9_�Xj���/��,?J�������yn}�s�)=��
��}#?l&@�(pHnD_e4��P�ܓ;=�v� U��o��R���)�����"���`���*���4���e�#�Vl%���g��)b�`ih��fovbJ�G>�o�e-��N}�<&���9����`��Y=%)�w�NYٽ����͗�*'�o�.ʣr�Y���X��J�=��������z��_�����A�wq`�d��q?t���3�i��M�cՁ��a�za�;qT�&
�������P��P���[]� �N���ᤶ��Ug�m����N(��R|6��7E���汰/0�i$�#p~�a�2��5c�I�l��	�'�*��p�� $���,���}�� w2�����{(�ݧ�^���%��ٻ� k�Bu4O#�3���4q�ɉ�"���	mEUw���wZ�V��-X���3Q�|s�нĤ�ޘȍTB��~��0u�ru�%�:�АV�#w-Ӕ�.%�b� �~lX���*��v"���^�~oѭA�u�0��I?�g1�b�ܩ��p�!o>v�͂$����2{{9?5�4\��4��Ė�<@���r�ef{��jK�
�%� >��1f��%�!���y�Da��5:E�J�hW�@�ڿ���[�ws���2z �(���B����ǣ-.�>�#_��T��ts�b	��=W����|����9��yo�/��BO]����Pl� ��M�zf�o���T�a��|n$��Z����wT��}���q2gL�9�:�˘hp�&O���e�����37$m�.#]�Td��MJf�����q`*�����[�K[���a����g(�A����6�L����k�������SVԪ���m�	6;�˲��r�Ů���-�r1-���۷t`N��z�����Q	���1"]nUUw�����eN��% ؗn��1PIg�eԗ[���א ��~gwwh]dG���ݥG��TU�x�����lD��7�X8��Y?�/&J�,������ק�,�̱ [���Hj�h}�����HH<�Wԃ��=��ny�_����ɛĴB<_�l?��K쟾��i�>_�}<�\@C���O*�� �W.&�Z�9.�h��'�8x_J��í�Ѵ���M�Dq�H�+�����<�*<�[��o�嗨��-bnpIT^*�T�S�7l�l��\���1����cA�o΅E�
����^R�NQБ����G��aS�ݞ�BO�&�n�dXŭL��;K�6T�'AEF�s����7I��1��Vfq�4�o��԰j<im"�E|D�N�Q����>�;F����-�@�Cm���vZ5�di}rc?/�t�����C�;�.�.�ь��ב�B1v��-k�0��;r5S��*Z6/=dh�N�NCV�/;v骗���@�W����k�T�4#dIƧ߹^�@�Rs��,�e/<7��5�4~	��#'�u��1�YÔR���4�1����
�L��z"B<K%%�k%G�:���q�d꼸ǁ�rX֜����CJ�iN�������FX��� �����	��I l�ߒ�����*9�[��
`���V%�}*���j:������8fF�D��@���>�aJ?!4>�r}R��{��-U8h�P�Ǆ�(�W�<⧕�d��8_	x�ԧ5����Hp1�Xv3E�
h�M��F�.y�>�z�WO]ww�OS���=��;&�8�����u�ubU��v'��{5�)�j�Y�#��q�<��h��q+oS�1������}�`�9<:�)fKr��l��6�&�x��7�	f�(-�WT�`����RU��tH��ɝ��ڒq�+�͸X�����s�>MM�jLhI^�L������2�5)�a@%��Di�zmt�h�8a0��rb��K��ݯz�b��)�=@2���vN�	���o��7�J&4�S�?��:2��%^�`�D����?*�队��@��V�xC��Ʉ�n��!�m�v��8W�kn���D���(���}"�{�k7�a;��ҥߤa,���6ra����i�Z���_�K���	����֞k�ıA�7����s��><�q�$��'��W�!F��oُϣ&��ט~h󸉨��쉀���4��#�����2\�����ߒke�����OY�H�iN��K��wj!Q����v��o-�Ǐ�bo1�+M�fT#�ԾzY�T0d8�N�џ�7^޷��6Q $��<Aftd�f�\�����U��o�S����eMA+ 	��w�}�2�Q&�.
(("l<VW��.�M�n~2����~�-�m:�%���@*Q.o���R�k�2����[��3�s�ʆ䢹b����G����:ۨ��"j��dq�S�o�w>Ĭ� )p�&}��Yw��^��|�*��Ԁݯw|X��0��9a+5oY��A�J�җy��4�r���{nY^�&�=�:���Jȷzs�U�9~1�t>�o�f�;y3�4���mu$o*��TN�J"ҿ�~zCd��0�8nq��=B��z���ְ��K�+�߼�D/D�d����1��}�H̚L�e��a�})��|Z5��b
�Y��#5(D�T�,枥���T��'e9ՠ���(���r�XlxVHYEB    fa00    18a0U�M�E�����T�
�A�N��nK~3#�]�u�#ђ)�[	w�qw�	��@q�?�6<m7}���Vf�ZF�����.P�=�O�o���Ŕo��~�Rj�g��U8�)=�.U�tEJ0�\�����(��{ԅ�6�u	���)}-�L�[���]�ڬ����EOX@�L�(��j^�j��*OU�G�c���Δ�z��j�^����/�.�G?i����<vRB�<�Y�䩋�J=��q�$�a�;�a�Rr	�óD2RSYe��hvn�'o��"����wv�b���q�~d��t�z]y�z��]W�߇�$�.L��[���C.�߆I�u���J�AS��67�"I�h�Y�Ry�P���s.t�1uA�-�o��۷2�������.b(��B�'�y%+�\F��]�$�h���MEw�I�{�1��r+�� X�/ꟊc�%8/ʠZ�]�i3��t#>W,�L��mȈ�'�Gk�מBZ�w���Ŏt��e¿�$�OLhf���ۈ�nH���u�C<v�'.�w�J�_��6�{Z�������^�F`yA�'�j᪢���B��o��W.��Jlm����~߮����Eh�z�b�<z0���a�w��{�-��	��oQ��F;M"�X׷�"G����}��gެ���M�i��G��s��I�vq��d)��(2�����/�Fnt� ����5��@��Ok��Bk���'�5<$��N!q簥9�П�9蓸Q��pkrj�[�L������]KwƵۿ��@�w��f�S���e��������z{�d���]�9���i=�ȼ%��:��=9�1x/������~��X����{�?�o5c8���i 9�y�0EO3Ҩ����[
Bt)���!g���DlZL��/���m��e ^ѝ�3�����Է~�u�8�!�x�c��mŲ��@s*6�ӕ�Re�;+-kK����p�.[+k��aFߣ
(M(#��j��"���u\AıLI�֪�}���9z�g���[��3Iߨ�����ʜ�=�>��N�-*�I�����=�e�es�Ae 3�lJ�d��d��' B+&L��m�����_������J�Ƒ.�^t��S�2U�CA��0Yq�Ŵ]�ʫ���s���� �8\_�D��&֔����&�~��KV5����L�	�V����3-uuk8�lN��s���X`=���zE	�4�,V���~����!YT�~�x\SK�)��N*��X۴cM��[h}�m\N ! ¾��_Q��ZV���\��|<���]`��dx��ZԐh��En��ʉ)0����K/�'��q�"��0�>"��^?@����x�a�C��9}�˩�!�1�+���5Ml��;ОJ&W�V��1�q4vr���d,�� ��A,�v���� �<}(~�9G�`�G�A] �������`��w�\^��ֳ ������M C�U�$>�bG�
ī�Kx��6m=�����f�d��W��*QJ�*m�� SE��W��v\M�3�I۩Z�l�^��izk�Q���?���>͂�sF��>�|<&��d���
����89諨��,�h��-�ۂ�?�B��1����BQ���C��ܵc�i|� ��e�.�0���nGyb�e�z���Ȳ�|���|Kc�f+��k)묾o�Bo\Gt5t	�!;Q��ʆ2&:� �Y��.�5���)uX�� ic���(�zT�t�.��U�n��2�Ά��v=��ә�"z��9ơio��µ�F"u�k�)[���N�f��P�P@�Gȑ ;6��食���d���〖����#���<B�hߖ
��T�{G]��`kT��� 9�w��B�V��R�!���Y`]�;@ȍ�·ƙy��w�ˡ�.r�F��3�(�a�@Q�eO�@?O8�U0;W� �;�1��jKҰ}܎ ��Mr�ſt/ߦ����J��h���Ȅv^��:�GlW0q�<��;P(���:�$���#me�{�C�M�D�&`���*?�XS[�͐Z���Y�׫�#�;��R���2*\�ׁR0��E��Va�6k������WM�(�^][]g0p��*����e���� �G���ڟ�����}Q�
��py@&���}e4T�-�)*}ۨ�'~4a+����&�v+S_�#L�*�Ȇ��˩�H�;ʵ��*������>�P�=2c�����o��j�����G���w��`��d��[�sv���28�U�_2�����Y��1<D0����>2�Ƥx2���n'��Ǘ���b�6�����ݖׄ����[Gv��h*΃Y��o3O�F�7G>)j���:Z��=��#)����k���6X\{!P�Z��6^��]�+��"�+�찃�9b��'�[Xފ(Q?�q���r�������6B�PKӘs�*�̉7'��Q�I6��^�>K����	3q��$I=��?&r04e�L�$��Kl�y�	p���{!�� `���M�2&�[�J"����4��`J�2=5�/[����$�CW�n�H|�Y���ϥ9�Q�ysdz��6ZS�m�Mbؿ�϶6v�,��a� ٛh#�2>�5�TP�c�{��Ǥ�U��(��tM�����9P�?�L.���R�N-���!e4*+���A;�Z��{�df#T�Ex�+�h㽻��d�y�Zǥ�;�K/�3+�R���Ԍ���� �*V�U�-2�	�<���=@
���ޜK�q��Nkē������ Ģ��-"ؤ�h&����@W����#,�pUƲ��VK�U�H�O��.U0,���j��8��������<�=|�k^��*�-��4IM��!{(��F�<��d�+�^v̞ÒE`<:?t�Z'ߣ�=d�h0�gF���b֦��Ie��H�V���fk���1���#�V:2q���H����MJ9k���iG4�0>ɒ�[� F#��玵�d&9�M�!{�t�Y ���a�h� ɤ���H_��ޙ�f�p�� ��})�̡��	?�W�R�nPn��Cw=�V��A�⻭H���$�Jԫ��2JŌ��O&?1O�e��or8��ů��^��c+v��/�wt���	U��n�:,��ǈ�R�$f�(�Ux^XAGi�Ak�⚾��3����.��Y���x�C��������D���*�'N��^��3~������X�*��б�2�/���|���z����:�	$Ƥ}��Fbx9'�򣊣D����h�\���,S��������Y����zel�ٶ{�,�?�h�_C�u ��"Y\1��+��<��������Jm��]�-_" 4������n��~Һ��5�r�9e\;�@��9�ˮ�Lj�$���A���<$^���!�:w��N���nb�x��Yrۯ ��l������v}�����e��d�2�lo�D�Z�
� �@ [j1>�(���¥hItqyl��j���|�'��T��� ���]0,��+5X�H[K��aKuc��*�Z�tL���>� �xSsy�> ]6�t7�?��������F�0O� A��S�T��d7ƂH�yΒ���E����t��l`b)�(!�7�KT�p�֔a�YP9�[es0^R���$��^O�h��
�����6+�4�Rb���6Q������\KxS���=;J��Ɗ����^=DfXA�:`�9�z�~������InI��x0���%�q��)E�ߘ��Pys-�-&6�j��UQ.u�d��=k���6`#�ܳ:ւʌ24��͒�9Ld{��B����R�g,�,f�]` >
��u�'�X��nS,DG�̾��- C��L���p��Y�����@��9��[h�?5&3��nb�b;nVs|�_��7����^r���1�_����7o���R�6������C�(PU��~�.�A�bHrWg���Ж�������Y	<U���}#�m�Xu���b$ )/�X���&��3>N���q�{��Vkz�]���o
8�4�l�7����D�l����
*,�����q����%�=;�Ɂg6��e�K����/����[F8&�gG��k���g�G<BIx��_J���>���gx��;P�*��[��0h�T��k�J���g}�Z��I-�>�a��t삈��2��#6��<�$"{��}@̣�U�N�P���{��������u{���7ɒ��wv�/I��|��s� ��ċS<ؕO#Az=Ob�y���4��N���i�$Q�:#N\������!=P���FP ��%�"�D�xԁ�U��ԯnb�<m��7	ޘq����9@GG�x\3�\R�r��´Yl��ӟ�������%,��=o�M�����b0��{�� �����4�4�.���q��l�׼�#$!y0�|���/��2���|�1$q�h�V�`v�y�LB�fod�����G�ԷX�@[���sP�|�/Z��,�"'�mI��.��k��Oѕ���:���T�ia��Z�ק�b��G!��yb�e��'�^e�1�����~�{���F��z��1O�A*�eN��9�P`ư��٬R}rO��X��/�6��%�䓸��P�^�w��v �Nv����-�^�*�BtUJ �@]����g��pc$Y�g�Ԏtk�1m�t�'����D��j�
8�)o@�E8v�e�'����G��*t�7�"���svvM����@�ڴ��	
�,�OL��2!�w#1%�5q�*��7Mo�/s9r���ҏG��d%?pcĚ?�uڅ����T�4��>ȇ���V�<�4�ā��$���U\v�UO/U�瓈���2C�9S�o�����&�:Q��[*�Ȑ3i��m�8,<H�:
%⻗7��4�Q�6�E=s�0m�9��)�LY4�|�3s�o��l/�Rh�S����2�e\w��~9�	U44�K!Ҝ��t�ůD���H�[��F��:�.���,z1�u����BY��
0?Np���V�'�����+�<�@���m����d���bk����{�ﰵ1H�Hzt��˓N��=��6�XV�]?�� ~-���j���ϔ�j�T�_�8��[Y;��Rp����� ƴ(���I�;l9g��qhb?.0ukK�ն�1'�Z�-�VMy��M�Nޜ��	flWԫ' �u���1ݒ�0��ɃD���y�;����U��y�dc��Ά˚}/9$�dԘ'��)�0��O��"�Á��=P◬\
}<��u*Q{V]��W�������y���nsB�=��L)JT�����Y��m/��!f���'�Z6�Y�D]�JN`�#|-+�!y�6�?Ip����i���d���K&J\p�>������� B0C�V��M[����������"f`��`��}
�˥�{�����IVa�`�W�=��V���b�w�'Uy l*P�M�}>�6&G(��E��X
S_�Mي���:�k�a���~+���_g�@L0x�e���P�G�oC}�8M���7������N���&?)U�d���)fӂp�m�a��h�(6�ۘ�9ڇ{��L��� �ae���z��f�	��s�Ӗ�lF��P��g�u6a L�cr�a�E��g��<�r�b�[`"O9@]��r�)WBA��t�)T}���T�>��^�hrn��ҾM���C�5h0�w��~�4ߋ-q:(qH��P���se7�)�z�h<w.(�w�<�)xb�����x�4�	��N?c����p��#��ׯ*�;����3��F��Yo�i�/��		˙�5rā��:�x�bma�X-����M�62��ϊoiC_7!?��$?���5L9Ł!���֯� �~Y���$8 `���6G����taط����C.O���
{���V	6�05K���ä�t�j�y�d�b�錮qF�L�I*	���&6!A4^�!��qS�`#r�y�(�ے����y~��X\{-qYx��G5��Lz���L�4g��g��&0҇_�R�r&&;���a <�iX�)W2�6�$ϗ*�<i��	M�l�+9�B�uSwf��A�h��*:^�j�4��\��ܨ��`��S�Ŝ�zy�R":O��7IcV���Fʍ���e��!XlxVHYEB    fa00    1200[4����#���3����އ�BG���:k����`�e��4���GVsx�VV`���q�O�QA��}K�Y�Du�_�#+|��P�f*��R��_Ӻ���n��-�5!<��)@��%�����nE���Z7:�_�.i�a�٧YɐQF�b�6	T�њԀ�8V���a��9�0���>���~Ps��E� ,!A��Y�e�G�R�O�����8M�~��}���_�hw��=n5x=�25X�hJߘ��ϓ� ���3����b�*��6iQ�:��]�e�e	-�+)�RZOWz��V V߯�l�ĴN�(����Z�b�����~Nb�!�[U�+A�J��^��U�sRD�W�f4�?���6P��X_���5��t�+ ��l{�>��ƻ^l�O�k�ȃb����Rg�0��d���Y2'�ai>��<�,��+�0p�[�O ��އ��ޔ�"e�&k��D��� 3: ���
���#�<�;�Z	R������Ѷ,�$���Ȯ��P���A�x�|S�>t��"d��4g�2�q�imY�0�2;�I[���.��8���e�=nf���\��	\��M|f����)�̀��&?>��+��^$7ZR���
�O��Ws4L�������e�G(E�NXR�d�BT=���1�f��%���කD���T�U�+Y9�1�56�Ȇw)͹���!���͞L����ڢ��8���Ň�^zb�®6�-7����I������W��Ͷ�J�t�CC��H�7��*"�-V���3�H�'��Y{���'��yO����H�JY�L`a�ٜ.�P�s/߰���ag���i}�I���&�4c�e�/�f��"���	�X�1"x���B+(��O�96�l������C�p�W|a�	 ��iN��p)~��K��J���ӯ}�e(����m��'�t_A}�NߥӜ�{��N�!PX����[��`t��~��Z��>���L�	8
&�;/G�U��6vGlȷ�/=�n/	,ef*:��@J�Sr5�)<���!�|h�cH}��z��U���� ��\i���1�	�v}���?^/��:'FJ����K�� ��$E��+�R�b���K�b_���Z���_�a��,��l(�!{���V�`��Qh
���e���b�U{:f�Ʒ�;J@I�%��������<�0��@,z�&��9�����b(sI�� !QB��
H3F`i�צ��A���5tpQf
,�������EA���w�!{�?�uOD]����I�E[>��N��/x�*�T�Fr!A�kVM��i2�2/	$�P�RM8��F½ţo�y��11ی�6;�JP8�9�C��td����x�V�髧W
"��������x�����W��ƥ���x�@���A����|9v�.�����ws�A*���oX���:�
 �y?F2r[@�|����}5�1�|�^ϊx��K�Ig �l�Iy\�;�ިq{K��$:4�/g�����<P�^bz]�=ehQ!��7L��'�7�Ԗ�)8�Z�-�,��D���U�C�!oJcȃo����QW�œ�H'-��B�iA�CicJ"7�ZP�r�{�Lp�9�L^��OC}1Q
�&k���Y�;��ff�rT��Muj���+�
̷#�$���rb�XL���J�
!� a�8�B�S��k���{��(��a��~��n_��f�ٹ�|���0�\��xJ�~��
$|OP�,�"�����u+>�<}|?xHd���.��L#]���v��R�.�i̖����c����=�?��*_8�+:�k��K8��~��a$0�FN��Ô�X�a��X���Gi���c�r��`ߤ�`Nv1�h�BG{�S�):!8h�����\��^�s��0lb�b~�D�����>%�^~�q�M��	���`��s�@?m�}�ɥg�ErL$3]��<�LB_������$��J��3lY_2��-{d��M-܀I��s? ���1<S�%�3��7��f%;�9_��٫�/��>_�IPn�����I"�	%��e;�3���^+1`B�y�(?����S�P�'��t2V�Y����t��Yp1�\q�$y.�Ua*rq]�a"���X���q�'9{@����F<ɴ$KlI�Q��ېil��[$$�\'$,���?�[h�O#��u'j�;?>&��k�:TF�j�O����~����e>[7Ĩ�(O�	���g|'����)Fa��N��W�y�[d�@#U�.�������5����b ���탚�g��?�276wO=�'˕��¡�C�b��bU�-��=��CuE���{`��Q��d��1�FFu����9��������0}I��P�%N�nY�1c؃,���υ|gY��1Q:>Z&K�'{u��PM���J��q�V��m*�ǈ�)�^HnIJ5
�cu8��u0p��<^���Wo�!I��V�_y|����K�������ng��������^�!�������T�\?���G��r4���:�D�Gc� �m�3uu�}�fV܇�,�Z������un��r� ���`�y��u�����~n�7O����pdOb���L��!=�)ó���>�5yl�j�v=���٫�K�j쌝�CsgM���f!�NP��nX6��"Ƃ���<�1�Uچ��[��b�j��h�[�"�ԛ'd�KN7���B�����O"�I�c8�h�Q02ՠ������? p ݿ p׸�[ !,��UŽ��l� ��u�iBPY�[>���Ż��ͽ1�nx�X8M���g�����t��>�,�Zד��ܚ��������i@�O`X|"��e2�v�;2�B�q��C�e7IE�&9�Ж$�`��K�j_P�4t �8��E��O~5�u��Ґ�D������8����>�y0�zQ��Y��.��l1���1v��*jmu�eb����_�wP4�]b�ׄk�������xI�SM&G�W�4eIe��E͘Q&J����2$dlܢ+��J���U��a�C��R`X:.���8�k��F�	��N�Q��`�6��� %Ұ�N>ҽ�W���Z�kQ���i�}���(�����*bs�n��P������ ��2odX!���Z�@�g��š�D}���~�-���WG���)�G��7������#.�%�b����:u�v���</(@^��_��fF���s`)�$	8����rU����|���ܞ6�OB��)���/g��᮶S�M��hf�V�ֹ�08)���@�+"(!����/OKP˩�0����um��;n���#�~E��3Q�!j�*氙ȶy�#3���̔r`���O*\���,��9�f��Qݪ:�3��o���d	������)DgTd:gִ�&���#"H�AÞ���^���x��q
�ri�_WM��s�4�#�p��%rcl��oDÐ��Y�����v@�m5i.�z�9f��ը�G;�5�{$�B!�E�j9i� ;]$?�7O��9X��i�Kr��F�����������&�q<�z}0.�$���B*��T�Z��ifOM�i�
 �1?���7��
����C���aRq�/�¾�,4�l��-7�@d�@8�Jx���|���l��u�F�i2Y�*��Ixp��˛�`�96�G�&a��oqz6��V��q��,+�/j2�o@���G%�P�7h���4uJs���LU�TGKM7�p�G�p�~�+��L䐼��7�jj�l�W�鰂�#А8	��켽Yu���B��(�`$\�`�n�&�t�T�}��#q�b�H� q����.2��C۰���F�3���R��f�3=V�|��p��D��N�o!�{��=�*��9Wؽ��(��"�(G��,��a��\��7\d��&ٝ�L���wa��nۊ��Ί�Z��F���/�^�i���I�S�l�Iޏ�ر�]��I ��Ϫ�����3�Rj� �5l�Ǟ ��Ab+[�"�r
��C������L�$����;�,��L�S�jTa���?�啧�i(��{�2rP��� �hc�P��s�zɵ�0�0��m�����Sb?��s���tC�]%d;�� $6����S�!������<�7����I_���@�
�4���,4��=D��Ϟz��-Z�/#�|5���g'�4�a�i�É�יa��9����;]/�L%�)
e���?0������+ ޑ���#${��W�M�AQ��K��# 3�Z�"%�-��˛�Z����/�� �[_m�p^)�2"I]�o�>f�{w_���(�3��` �kTp��{�K��Az�z��[�'��;S������z
.BjB;���OW�H�m��Mc�[ ��I�'Ɏ��>
u?���@�����[CE�	�觀6A�r�A�=�kő��a���uڅ��S��H�y,?F�
3�[z�g�V�s0~b�(�[�~��a�Ƹ�5�vl_Q�ʈ�|�yB��5��|�����D�֫x|hK�ʇ�X�bphXlxVHYEB    88c9     8f0�9�d7n��*�7d�i� ��hk�T�hi�U�KY>��8�.���/�?s������u���Ǘ�'n�o�d��`)hma�a�� X�u����s��}W���w�I\m�8I �H�R���N.��FS�!��;G�P����(�xB	!������*�n�.'�7L��EЈ�ۤ��2驺f�ti�>��sК�veU��5�d6#O���fd�%��!���tKd��vD<�݌�G��00������^��񻼍��F���9͑!E�}N��v���QŔc��U^�f� �
k�A��a�w5d/A��g���=��Fh��-��]�{ d!���%�fwK�/�.buQo�^y�� �푧�:-�&gLP�ҰMnJ�+lx� �v��&]G3�)��Hd����`̈́J�J<�]s�i���f}��\�3;���S�
p�����d�y����P˧�������65vկ�<�+����>"�w����z(��o���*l��
^nKd�}I%:�Lh�ө��\�xt.���k���ٳ��O���V��3$�gk��:�;�;3�Ը�F��`��C�K=��?�k0�/ri�B�!Ӓ�,-U�#�́����ٗ�*`Z����3��JY�x��D����l��"%�V\M.,��$6�niү_H~#(�Iѽ�#�����Pۊ���m����R��f�B2�����=�O��(�Ř��2L\SAX$Ɖ~_&��El�Z�i��:D�����v�0�@->����&N5#�Or��O" 5���%;a��8ϣ����To��.Q�����괁4����T��%�&��7��Ƈ����G�Y:j��V`_�Ӹ.�WD�$~E{mOG9?�5�[A�x�jRd��av������RT�&5	B��{U�Y� �%/zٔ?[�)�ڸ�dU�a�[W0�'����S�[b�/Ԍ�*���g�d(s�r(�|o���2=N%����@:F�Y/��&��#�eM�S�e��Kdj>�!�|���X8�@��q)�)�
�H��o�#V�s�C�NN��5s�;�c�<��A��_� 6=}��T�Z�gA�r�[!&��$M���k��UI��!�z�|�c����G<8u~zq�Tu���x�c��L��@b��������wV�Y�ĳI�ؖdw�dڟ�N�5�&z�3{T�Y��j�n�� H���,� U�Y8���jo���4Z�Fw�*�aʬ�E8] U���=����F=�}|==�qtG��'�-�?ƀ�Ӵr��d��w�}g5q�po��D�䐾��7ӿ���C՜cW���u��{��ֽ�S��� ����"�r�m=S�9�5��4b��f�!]�t��"@��F���[�K^�����H��mؚcl�.�.㢍���2YR���+����uKm��bb	��Av��(91�����#��i�T���އ���*�F�K�YҜ�9#���ސ�ՉK�j�N��d���ϐD�ŴZ���M���v�Ɩ�v�1N6�,�O�y�^agv;�V��Z�%���V���
��=}��V�i)�r����dsg�03�:��!�q�6 �������S�"��sO.mf���9���q�j��ʻmR��?\�]�b������Az�W�C�?qC�:�[�>7#����{�>x�Eg�� g7~��=���b��Z�T	�$D��jgn=��W}9C~}�z�[�7�#�4>/m���&i�n�CQ��Lsx��J�D�)�\a��w�`Ҷ���1:�ƀw�[m�gg{��'-6�:���:��>��f�s�0ηp��+w0�TS����o�|��*�1�%���p\#"֑��!xr�}x@��Sӄۜ��?V����$U��?@��֐W�Y�c�q�� �-n]�*�m`tJ���>�E"�x��?��Dj.Җ���i�2�BN5 F/���|'����W��B!����f��|EM�w�� ����~�ܧR.�&d7�IM���Ow,UIK�6($pB��Bz<�͈�fv~���D�9�ٳ�B|�U:C�-o(�V�=�m./j&!v��P`a��2�(���y�:���/���I�\P		�z��[�6��D��_��a�X9�^��u�3��}Iρ�D����DkN�@��9�'�Q)�\�_F�l�x�E9$�B���.&�w���.Ԩ/a�I�9g�j;�#�礬� �`��%�TS�ié�Κ����zc�bc��Y�,�\p>