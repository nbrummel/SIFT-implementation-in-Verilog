XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ͷW��y��yg���A���}��*|���\1QM_��m4ϧ]n���x���`>�$�XB��l�ݫ�r6�O'?72�9������=3*��r�@�̤���DF��m����%���9��"Lqyd���6I�}?��.Ww_��[�� �/AOG���}� ��B�YH/�?� /bsv�w6_̧��ǡޜ%���ms"�$����g�����:��K��=��s�&�N8Kq\
z���>���qXM@z*q�A,'�O��v����W��6���S����]�_о(u�vM�BX������]�ˀ������DjFGm�F�/СW��9i�{Ӹ"�����z��h�/��>D`Ľ.�9��D��@c"n�r���\M"�,�#WqI�r�W��D`C[u�@9��d���>J�a�>�xC�n�B%��1TW�T���d���-�\�(��O��[q���H^��A/d��V�t�g1b3����!"���sÎ�>�:���������W�5���S״"�������jzQ���tv=����w\D�'&Qp�xGn��2 ����=���/�����j��uD24M���!o�lLݢ)����`�+��UӢ}f`#_D��@��>���"��M�6�<�_��V���
A)��p:�vV����1%�A�1�;�'�"eY�B���+	ؘ�(!KNqf'Ok�`9���ғ��)�����jv��[�^t�WZE�PP��p��3�WuXlxVHYEB    3504     cb0S���$��?�[�ϻ ����)��<��J�7D�I�&�Y?�\<��yR�u�%�u��a���1@�ߌ��j��s�Sq�r�Zc����9e����9�3�mb�X�����AMƞ���V�h|'I��W"}�
ˁ��E��/�k���mm30�P���M�H֋DT��V[���9o��ʲIlM�eb�C�X���� �	���V�, �!��L>�xg��Y���+<L�L$�V�ǹ�`�qw�k���Α)M� ɀ�a.���s��~�v��_;���-����_/�9`$�`80g�p�������	���R�\b#𚏙b���$OGre�NM���@�g�#9H[�o`5��m��d�7cct\S2T�YԻ4�U?�涪�?����G�#7|y֬�ENg�90�n�DV���G�,ۭ+�ib'�V�y�� )�)(�ni�^y���=�7o[Ř���%5��$�h�}2��2Q.� ���;�6�3燉dx�a���h�Ì����}ￍ�1�j�#g碧	iG� R&\źP�$�E��]����ƛ�,�D *���<�Bw�;M�R):�#�Y�O�U�I�6ԏ���R����Z��3IU��ԗ�-^��p�b��� 
�f^E��i��p+�
U��J��'?3&�Rw��h��D�!�uO�FN���*lV*:C��m�����Z��x�>UiSh����r%qkI�\�x�.�J|*�Np�4��sB]Éw�A�'
fH�[���_#~������I*���fl�k�>��z�Ъ�v���4D�9��Ys�e������:?B�/��-�d�OQ�t�S���]�1�c�uMd��PlPy}Q����N&P}��r�\�GO������1�y'�c�Ex��T�WF-%{���*Ed&8O؍�Ԓ�y����8��[�%lɎ�b���{�|T��F�U��.���Vd�x��B��?O>L��
������'9=�#�R��i��|�3v��t�*�/�+�w�:�Y�<�h��>�]S�*�F�vӭ�F��4��j�A�qm`P��vYp�=.��1���m���Q|s��|1YHa�ug{]���&)�7E�嘷[}�b�4^P�����p{��ٸt]�n��$U<&ड़�gm�?o��m����Gq��j��T����M+o �Д��Sr���U�����������l v�%Q�j����I$����&w�Nհ��Pc�]h���^C��9�� c��$!���!Ts9370��#B�H����$U��Mz��&�|L����<|�}�:pf_	��2#���U�%��Dm[F�t}!0�brA���M_UM��mȈ~cUĎGY�M������`��g�sK�P�j'��.�fm�I_�o����P�I�n��ز�1�"�W� �ޞk����?�l�-��$�2����2o>ji��0����t\��P��MmY wd��ˍ4�&2y��Z�������Y$'�t6v�l�030�UQPKibs	i�G�v��J�L]��MWy%rp�	D�[��D��x����¹�$h_�x5K	�����̕�e"]̝z�Y��b8��*w����7H���嬗�ً��V[��A�qA�W��_S�8bP3�$OdZ����<�(�EOz����6j�\� �Op6Y?r����N��$\�$#&L�tgҌ��C�{0���;�7���b{���F|�|C��៕�4�b8S��b 2��B�|���3��6\� ��O^4W�����@b�e����X�4�jӯx��Gُ�U��)���0���ҀK\��*���c>���I�r�l!�1�>��Jo���%�J�Q�Fٯ�s���Y�����8����n�v$k~���_�`rx��)����HC��Ȇ�	4m�|q�Tw�Y��&�K-/'Ȕ�1�u�+sy��k��)�V4[rv�q�9i#�\���!r��  ���ǯ$�/!���]���j�D`�{��J�w(O21ПBYA}i�u������u�VG݃�):����e&�sKj�z�2�pc�6%><Mh�Z���
y@/8�-�#X�Y�G� }N����W��-_�X�'�	x���t�1�pb��xg�>�j�َ�f6�n�k�՗	�t�?)��#��=h�Zϓ�m�� j���ZF7����2���o��̘�|�BC�d�-�,j�0^��ՔM�<J��hzi̟ۺ	�ǫ�*h�����9'���,�i���m^! �J_P���ߪג����V���T��gH�tk����pɐDg����sU�7�ȡ���'R^�Y�h�85Y��*3`�a�j&�~ᛩ�h����W$.OT:��+Y�z��P��1I�����Q�l`M9�A8�q��\`��`��͢{Q�B��� edz� �p��|+�l0&�#�7�S�.f|�Ӷ#���e�É��m������Yrz�2�R�؃������ с�g�����Ժ�� ��.@�9�+��a9�Y=;�������p i��`���
��s��_9%/���l�!H��4.M%}(���לW��y .�N��������I��w3�$�%�Yʶ�#8����s�0��#�=uy��N��=Ndo1�^r�/kI�qTrl����0W�2��{�ב^8�ZD��� 
{�0Bپ$�ߌ}��5bX 83Xv36��5�~P��a(����nxz�q~*���k�\θ3
�x%V���d��U>(�����͝��%�P +�5Y���
8ޙ���a`{/!�b�}���1O������v׸�r	9�O�"4��&�W�C=B0r:Zش ^� 2K��\.46�=*�][�C1os�#t_2���������0ߐ{ľLe�L_ua���)>��#����b>�򛜇@Y�m!�!�C"P#�s.K}�˄��;�n�@�$�0�׎�(mkvR�op���(�=�e���M���>�/���2�Y���'�)� ���Ӭ-V&/$�X�d�ߞo��3B���gӹ�.��5�D��/�S�d��m��*w��0t���PDP�C]���7yQ&{k���՜V��@V�T�%l�j[�(N�?1?�d}�O:"J$�'���@�Bxۭha�<!��81�y�p"Yk�0ۺ�G���˫��b|h�HP�橝�7�D4�� #hN��Hc�}l��>N� �x����7ϝ