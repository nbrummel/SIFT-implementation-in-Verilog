XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���U��fD���H��w>U>)�3�|b_��
8�W�n�dre�g�e�d@��~a��4��-!��I��K\�FU���5�Jͭ
�&�,O��h �ǋ ωS�	���
g1� h`5꾉� .��6�!���ۚ�K�� G&��K�������d�,�u�ݵ�o�-�_��y����:��=CW��*��fϞ���eC1�e�J��P���E/���~��/5�E�&�R� j)�����`8IYBF\�~�������L�2#+X�0+rZ������Eh�� 5ְ$SD�;�=�8�Y����gYB5�į��n{徢��Ş��ne��T\����l����a�n!�)u�U#5���&�� k��s(�u�s����,X&�=��������C���4�����e�Ҁ�/���Y�xN�9�����y<A�s[N����
Й�T=����lmW^|'@��
{�w?8�ϩ=,4؎�g��=ѐ��E;�z�چY1�RmF%�A@�ߒ�=�w�G&�l!�+O�%�T|��~,�?�
�n��!)#��2AJ<�sEi*�A;�40D�Q�#�c���U��#1-,�$�)�j/z]�_�|��˂UM0�1/�*��a�}��4
����sك�*0����ˣ�Z�k}��׺8Ě�1` 2�ϸ�3��M?Kb�F�TD����ݷp���I��(91h�"))M�B*S7�o*��#ր�k	)�̢�h-Cϱ�G�QܹUm16�ӓ,D�TKuf�XlxVHYEB    4192     dd08��n�1I�+]��1bd��#˓�0�<~�)"�k�y\l�9�Q��i*A�O�{�|6u����̶��\�� @�W毇N��"��`o���d�DA�8��5"/���	��ۈ)��YFbMĩ�	A�6� ���P��
����|��7��'ŶP�t����_�kM�����Iƃh��v��mi��0Phk�T�y�PG�\�c���5�g��P_z>�l=NBy��و���j�w���>���~�f;�gQ��t�_ý/����= `iT>}��K2vE	�z�"2W�ڨ<۸�2�%�Kt�,�At�I���TA��m��C.m�2�:e`4ß�X�m��LL-�YT�H���2*r� o��V�w����S[Is��dBd�Dv2&�xu�o�L��"c���Y�Afs�I�bvl�����ijt�a9���Q��b��#�"�m�yvpLX�iK��w��䬃]:������99�\�-�Bͳ�m��4v�sAD1A�) �w�7�n&��ҹ��g���桞v��Z�����>ګ�ĨW��?�bP��XX{�d�8�R��}~�	J��4L�&��їY��It�-{�0l����[�XO@�?��A����G�j�:��quWPUz�Z���h��P�غ|�4Uae8�9��DW(�����$ND1�^�uj��ED�e��,@6f�ƿY`�N�[8��6�U�4�����1���#"S��K����xU6����p��r� �=�j�x^o�;%fQ�1��)��}��I-sAa������z�-	�����@{�	%^����17��A�(��h��΄s	�=�f/T)�H�	&
����E8E#�����)v�+
��f}vs<��d���{ӧ}Ԁ�{�7� ���e�Z��T��3�R�E�o���+�j;��a�SX�M�3Ld;"�A���kƘ�9X�� ��V����9�� ���dE��Bg,��S��:iO�����ݗl}�������i������Z��va&��톽Y���IpLc$p�c�T�I�$��'Z�n�#�{��G�*�N\~b/s�R�(������!���л:DQQ�=�4�s�/���5s��j����9�VF�j
e���ή���_�ܖ�6>4wd
y�����tx=&9���B���&A�D�m�C|T��3�4�݆��-��D�����`M��܏��HB�����7�ɷ2�,X%3����W�F����B�`�yP*��'-�C$s�0d�47�>��M����7���nF_��J�GA�j�gY��΢����C�WT�T��|9;:��m:i�������ԇ���4S ��ݳ�l"�#z���a��� �����9�)dݟj󬌖�������Iݭ-��cO���ݺGb#oΡG��?���_ɳ��dK�J��`4���~U���n���QH�Z9	��g:n�
��������a�UbAS]�SU��Ҙ��{mv�j��}F��y$f�uK���*nw&�W7�}� �^Z�t"xQ�
��t��н�sr�eK�w-����� �:z�Rc�H~[lr-� �D�genh�&�u����g.���	��PGa�%k�U!7���U��U~b�]��ib%�&�9T���6d���,R����S�mT����z;������O5�h�����n
k���bێ&u�K_U��F���yYwS�O"��ϧ!�R�`8s�w��T�	.T�ڻE�0��⳨��٣G=�B��/qp��ٺx}ێ=}	~x%�z�;'=��:����#4��6G/�u��y�<KJ`�	w*�"m����b�_�)ﬔ]<|�����Xƭ��[ZF�ܬ�(|K���ꔠ�H�+��BQf��B8,�O�o��qL�g�P��V.�]��b���I� �~�{8���O���<I]�?� E��K7`J�~Q2��w�9��ǍuW!gd�&��¬;���7�T������;˯�rNc��P+��'�3Й*�<3�)�����ƀ��� ��&�#pm9�ڻ�鐜�'�9BE~�P��41m/�G��9�e�؛�w ݈����~��FƄ|ɣs��-�ۮdO�5 '$���`�w��y�k�L��k�����֎��`������lI�J�Xr��,���J�\Y&�W�;�ƶv��6�T�PqU�N�Y��[T����&`[v�A%�J�uJQ���cq���� H�X�{Q��Ek��%$�*�/}���c��(�:�*�!��K��++6E��������������Ǌզ��1h�:卮Nަ��GIYn��Ӧ;�#OA;����C<���ι�LИ������jn�1�����\��]�d	q�B~X�8\su�~EDpR_N�À�BE{�z�_�[4.����=���m#���FM_IY���;neŵ����Ys
�4�g�i�=}A�q��e�9��f����:�*�\�R�����H"�]>WWB��G?��;2��T9��Z���b$�	M������DX�M�!��_�pZ��` ��'�c���!���|�k������>
3v9S�	�X*n0QV�4�ՑuZ�r�T7z��3�����؍��@�0�pw�q�S�LmQ�cX�����6~'k��E�$�dϟQ.ǍS�k]�w��(��G��������~Ɩ^�L��zZ%+��ǒ+Me�y3���G�R�t�[mk&d}t�H!̎�=ߪ�4A�>��?n(KA��������uu�|��0{��^�}�;�e&4��]������6AU�l��
x��	�A��P9?{�q˨�ԂO9�K��,,]����b�(�zw�F����-}�����}�
�ŮU��j�,Y��j���e;eh;�ǥ6=WWL.�q�C�p�x�����R�*~�zW8�q�dƏ^#��\����դ=j���nG ���c��S�-b�;T���ϔk�r��"b�$*�y�������Y+���ӱ'u��#s8:m��i�W䊘�v����9���maa��+�Z�lTJ��_@]�����?!�舰�>E��e�.b6����k�a�3�t)"8�%#_K�|WC�l9�h8�m�R�Y�QY�MP(9�˵l���Y?����Cݝ%u�^��\8�o�z���W	��
�g�G`�Rby5j�4��S��}:�%����(j��wZ����N�"A�5i5�H&`@EH��'����ё���\��, �kBy��z�>����{�dx���y�M��LM�kb�ff��6}@�M�
U���C�Eq��]�K�9�@g6Z�j��:ۤٸ�'K>n�R�� 6^eƈ�ZR���W|���ȤF�{?�>+[��Xx>h�9Ü�a!g�?&��?������׭ߕ,5i����"V�.�@U2�%����f�۰����	O��^o����c)`�ծ�Ko�	�0�3&���a�
��*�f�
��i-�t$�]GU!�Fy�9ix���_G��Q