XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9�FMuGm����6v�Q�8�X����"�_�?�w?٪4�*:	=aW�ݡ&Z}��D9i��!3�!�z��8Ɉt,�����*tP�&�m��7
k�+V���#���H���`��,|�J E���8(�p�X�c���#��d�|��+���-���+zyYދ�C��VP�	+�{A��-.���W,c?ܸ˺��
�j�G�ODi����i������҅z�0.Ə�'g�ih�Eh�%Ao�4���[��y�Ew˫�A5�6��?�ȱ���,N�����]�6U����.$�ȧsĉ��~FX)0_E�0���gA���%ח5�=���MC_2�xƷ`j�U����U.�+�a�F��0��W �����-8Ppn��'$��ɤ!�	;�_��s�>|�j~�WHxiR��xHe�،����I���2S��;���iM~e���8e�T0e/�V��j^ƛ��o��;u�2ƚ���J{Ɲ�� )_d*��:4 
Α��)��O&1F>Z��k$������LhC�Y�壞���I���������R���`^��)1X#�� %z�N��r3�@�;�@�?̲3�+3ޅ�+A��	Q���çY���9}�B`��;��Bt^�������):�K[m�9��j�ϋ k�Q}�	�5��R*�
d�䊐���"c"�+u<�`X �4	G!z	jd��J�����R�����О�xأ�Z݆˺�_������U�s&��XlxVHYEB    6cf0    1960��Px#MV���j	':��NWTH�iU����8�dh
f�o]%p�&97X��a?�)dK\wgGG�����uyR���QjG�a����>�+9ޘ	��i�	�
LyC�)�M�!��A�1Afi�����XgK(tQ�H��1�0��I������dn�{�)V͒��f��)*WP�GL�<��;R��Xcȇ��PV,;��9���y����"p�K�<���SQ�����Ω��Ai�
�ݾ뵎�秕�XW����4Z���v� B�Gs�'	��U��Fj��A-�L���,XW'��I�Y0��a�|t�ֹwYZb2kk�:L���:���|���D�H�����"`��U��dBj�?Zs&��X��Q��H$��]mm����ŗ�/�z�jPed�����w4���Jpn���y�� NY��0���7���4�C�!zvk��ظr6���M��������C��8���LqLZɖS�y��0�L4��%�.�����fX8�9��a��f�>�\��L��ʳ֌ޗ���΁,]F�C�f=������m���o���||$�X�/���+�)7�S'�j��Αm#��F��]��o�տiDO�D�����Q 
�	 ���y�* ��D� 1*	i���<Kt��d�L��/�4�nڑ��8�t��Y��+�\e�3�e�E��>7T�Ӣ�a�1p�XV��ρ\�w\jH��H���c4)��r���1�r�Y����ɮX��-:#-�`e�n�`�qi�?�\���g�ު�=�s�L����y�QM���x�{�A6����\���z��j��׉Gϩps1};����c��I��:Db��TΊ��{V�3�`l�F��N��۳��vO@9�;^��^�Gb5���4^�<�X���e�5;�9nw��
e�	�V�%�w��w�\N~�9B:�Ea���a�H�41�۶Ʋ�3>�@�2w�b�2�R��b/��D&,ЗJ�C��C��a�u��gݒ.� ������V�ĄZ�zfh;�)JPXA@�Fe����`e��n�{���׊z��Ã�%�e-m��Ƌ�**�R����,�p�99*�_�]���ΛF<�*ʈt�д,y��U��O��:RF����%���5��r۪JP���.�`{h���tr����s�V=wgF�8��y�fs8f`�S)���w[WK�UR���M_���u؉B�"N��M�0���.q����T!��__�n3*&	�`��w��,�Z�J�9A����m��"��p�櫾s70��r���{�y����&�$��I���\(��,i�ƪ�J[�����E�r��s��#��n(���T���Q#f)��?���U�]h<������Li�q?�]Ns��?17�f�����/��%=Q�U���"��T����^��]�˃y���8:���^���2WE�P���x���"mpT�g�kK%�(���?%�ě�.!��C5�؁�t.��t��U�=�?oX2Ԝ���4���J�0~p=�tf���D���Gi��Vr��d	6�r��O����h,�;�v�ח�&|Y�� ����y"��8m�þ�&f�B$�mk) �yQ�'�;�d*G~Y�-��W�s�}�S^;n�����㧀.�z�:��Nh�& 2w;�,�}?tgc�/��[�����pXJ��46i4�g����'H�8��sOYhi�q��I��:��n)�)���¿a���!��Jl׵g�0k>k��E{8����0�K�PT)^�3N~a�)��c����?�O�gј�fb�捁9���-L|�{C�G�;�{d�)*"9���F����Td<e�I�8!F��p�)�g�)�V�������5$jS��S��\^p��ԫ��Vt_��c�a��"\:���iv��B�{L�J����};TX�ޜ�vPdET�2rS��k*#>I�˰12N�%��C]d�9�'-�3hqE�ߩ0	؎��yͪIɓ"���X<��&��Xdyk�ѫY96׮���T>���\8��B����In&ݓ������ T����`qE}A����h�����=�?KȈ��MîN�'C����|2�sb �[�s��a;G�(�,zY�Q��u �~�I�L4�ύ=�Zf�:E>��.kYt]|'t.��n޶b�ܠ1���,A��s�;���˾��P'
��ɘa��̠�I�xukx�A@o4lC_��ga2j7bhS.�G0�����q4�������FxH��IPl5N ˠ�>�@l�Q0�8GWry�C�ma�d�
�F��u�?\�p%��{���6cE.�I���^l��_�֍�-:��3���4ጮ���a*VZV�������vZj��� �N�d�����ײ[V�(����f#+�5�٥�E� l�֝�X���Y���n��0I��&Go�;�LND�3����o�S3�$Ġ�C���u���2���&d��A��MPv�Oԃ��=�zU������~RSW�T�p�'3DK�A�G�O���f�-L�{P|mx^	Ɠvdʙ�P*�7��Ct�rb�(~�ĭE���hO�_��h�PkRT��_y�z~=�� �����HCHO�������W��>�3�(�m�	�|�n�
�]Ƞ����oI�B�Q����?)�Q��* ���KSRA�:r���f�h�}�Y\�Ą�Pt����@��s�㳿�g� ���rE̐��辂C�(��	e)QAީ&(����d&^��%H��d��Bʭ������p#f���� �o=ѝ�	½\o�b�`���+��zj�x�!^i���ަ����̉��{Nf���{a'��\0w�'D�9C�'�TS
��,.ˉz�@�Y�����F^�}�k�^GQ�ژZh�빖v�q\�B���/S����i�2�J�4�x�
n>�d�;�]%��ѝ��wsa�9l��p�.��x�*T��98i���2����9^VW��q7ƿ�w�����F�)s7K'2�-��C��
~�;�	3=�]w��� �I�K�4q�t�&���f�<+�����/�a-S����㯊����չ�J��J�].�L���ݼ�x����Gw�@�ޮάg�0�a��	#� EPG���d%�U��P.([���/פȭ�Z:F�0�i�
Ee"��(��:3�E(��NZ�0�պ�g���3��)Ċ�@	��̄�AMk�j��ś��-�eaM/����&�*k�`��ć����ê~x�Bd��+{5����{\�=)��6����Cc�_�,�Sa�w|V���|�sϔO�D�a��^��K��i�}�c��pS���ҌG�4�D2�i��\-W��h�2ϣ��w;�[c�C�_�&z]n��q���nʊ���m�KaS"�	��@k�ݛPt{��@�\�8��,7m��
Y4[���R
9b6WA�,�7�%���蜄��.ZM�v�;��ZlF�Q��wh��Y�������:t�tޝ��|P�~l�N�C�̛����&r��x��C�6�3�g�ND�a2���N�� .�U�ݫ2s'�<��:���2��kdHV��! �l�جM��v������6��B�ez ��5b��s��`�Ñg�L��~��1�8W<t,���`LT�|롅���F=R���Ǫ����E}L8��G@�K�l����O&Z ��jYz�\�dRۻ#=�4t�k�XuA7�ީ���C�f���,��3�{'�(�qr]���ۭP��.B�N[��7�����ݠ=�9��އm����Ԛ�1�XP��j�Fw߾�EϤۼ1
c��\�]l1x^$�x������L������pҬ�x�Li�=l�K(�U4ڎW6%��8�z9��{m$��$ØV�Y�`�!_O�o*�a�=y�1iU:}���.m�h:�5l��@ejzc���Ч���'����T��qT\ l!7�>�V��A(�,���۞ �_~����ʟ_��C��� ڔƵ�P[���ފP�=�������Q���J!nbw�G,X`M?,O�hJ|�׳��x�Uj%`/�&�M�{B0�V���������gs��J��:*fZ�|���L�ؔ�h^m+���MBv���P� �����E�%ә�Lձ��;���n�"�;8�X�	��2�y�Ӵ ��2��'�򬣬#�W����
�`����c��B���V����^`�ᄶ�'V�o��u�*�:����;��0}z[���p�'hr���&��\UW���gk���LJi_ I����Dn,(�Z&o�n�	�lI�2�!�BI{�Qﾡoc���`���)k&�7��x��4A��2�N�`m����0	� �k=��Qt��irim�v 0���zŶ�N�;���g��JV���=3��bt��Zl�'��`�pċ�[Q�=�zG <Lj�P�	��j(��Z�Q�\��Jg%�'��5�q\�_y���p����"R�:LZ�y|q��Z�D�F��֭`n��~���.`\�䤾�ڲ�A+�����(��������D�-������t�
��DR�Q?�g�0,S~�����fq��|[�r��ywdt�����/;,O�����q��7�t~�|TR�\�l�O�z"E\����<B-&�:�)L���$8�<U$�ۿx�Yg�b �뵣����ӾE�К�>�)�"�x!9�ar�|'�E�Dl�`^�g�\2�L���}��]�-ݺ�N����-���n/"m,��/�%����t�]k�8,}Oѓd�� ��7��H4��>a�˞r��l�m<�ڊ�G��o4م�:��їh��2���¥�)��V�@i�.է]��0�Q��W~�̟���w��%���F�j�S���.-�����o��w��N��hk�=3���+��&<�X�泤}�N&�l�-�����_��OwnU����D	��",�m7K}�M��Ez�M���yֽ}�B%��e޺��C�(d�XP�<�v����	"��,�M�-1�0J�1^D����"�(�'á�xl��fi�&z�Z��9p���pBJb䗊d�{g9��*q;�ر���Ҿ��y	QYR0�(�~M%U��+�I��P�tq����T-���հbj��p��o�@������J<[���h��T�!!%������O~ج���J^�}E<��9���"���:��η���T����(pe�QM?��(SN���[�OO�Z���N�b��"@^�oG*h�J�y~2~��VA{�y�\5l�P)�z =4�%��EC@?YhJɧ1�}� �x�Ge�65g�m���L�y]�X���G�n����������jtY�5BI��r�����+���-^����Y����������"��Uyo�[�(�[�g��`;UI��� ��c��$�-��:H��(��1ݮ������9*�3����Vx9������)�ߺ]lv�'�������}����Њ��7��|���{����/XAg��'}��.7{�L��8��@������L�"��5|E^�!�=�7X��:�m�������U{��o��bɦ��n+8����TsxI�|u����x�Z~�N�BL-

֕OA�Zj�ZϿ���&�;F����B=����yNPr�c^�^ȣnI�n��T�����rn5 +Ų?�`����,em�����y]" 6=]�r�<P�ŐU7�i�ρi�V��b�T�:���z�?������|O2c��s������氄�M"���J�Ϲ�_�6Y�;'5X�Y9�u�ӯ��%���Y�~�N��X��Rvx�Cng�����n�B��c(�	n�����l��c/��x�)k�gj�c���|`DZ!�SY <�Q�"h��l!]�����q�A{� /Ҥ�č2���e�`� ]R��>���
=��{����m�8�����#�"�o�{l�r�;���)V��{���n���W�4��$t>c a4ht�6����@Ϊ�^�?F������_�l�H�}�S �:ǂr�j+����E<OÉ�1�`�y-v�@��J1��u��N�tNc�e�<ç�`n��,��b��2>���	�����F�;m�c���B5:�l�}i�
;����ݟopZu�[���Ar���#g�̟�J3ȵ�7��*���zW�z�U��(t�,?�J�(V��%�c
,�(OIӽG����QA�����l��^A�u�KYS�\K@9��1�fQ���9��O%�� 2:F<Z��Uq{��hʜ�����F�D�*F��y�L����,�n�p$��&��;8�Oyt�Q�g�D?��t?h�JH�S
й� yv\�u�2;�.��F���I闉�M��>�@�`��2Χ*��