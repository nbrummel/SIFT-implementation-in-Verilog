XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��# �6iI@!�������y*�0\�yH��L��e廐~Ж	꩔��˓�ߠ�7�!5��l.X%�����(��_`��$�B?H��x��%�s��ww liw�{��5�ݐ$�>���8lB EsU�Κm���ԇ����bg!�I�8��Ɂ�3~��TI'`h����HW. Wd\�y|�5��G�l�}�G�mQu�O׶*{6�B6�dB �j�'��JQ��Zݳ����Ai1�a��o�	T@����o�*^>�����~������������H���):��\�o�D�E�4�j����(^�&k#�7�Ř�ޑD$����#�
&Z�����Sy]�\�`A`�Q�F�ڈƀ��J��K$�%~��	����k��9L��-����\&�6_�V`ܵ����HD+G��uq>n�";W�/���R���F�� s��'�����af������*�<`�(�8�s��
���M���>Ko�wk4��)��-�[0c�ˆ�v�s�d�[�4h.'bɫj�x�Lk�!��F���TT�-��=�*�؊�Y�+��1���*ɩ�s���I���r��_5�|@C��f�*Jw��^�u�Xm�%0�`���VB�Y3BF�������#erA�e[@X�V%n��a.[9IA��	�xTrpJ�C.�7��RQ��2��:"kmH�E�*\l"Ǩ���jȓTx��(��Sⱪx��\MP(���A���������S]���6U��R?��	\8����!��XlxVHYEB    5dd9    1240�1G��ڽ��ۤ��Rm�`Z�fKTlpe7儠Nl�h56:�A��)(@���v��"��f[q��~A�t�hE��i�m|�&a��u�$�����!qİ~��{j�+���d�PS\X�(|��R��܋R����|���ח��W��W��L�tIF������:f�i$X"4�Zޘ�M4���4W�����iKF��Pc\�SWY��%�,,�	��k���B�ՃC��$,��h�F�d�:�4��a��n��q��a��_5<q��\��q��?�Ӱ��A�H�|��=���z����%� �S9�J�њ���Kޏ*�{X��T��bi[B�,���Ű��V�����%�h���^�mF%��e*8����Y\�7�Y�d��M/�H.Z:�iE��I�cL���-�.�0���?(�3�H�O�=綱ekU=�ۊQ���� ����Tx!�IS`�:	�qB��!r΍�E�b �+Ƀ���(き�uH>n���������$�.���[am ܼp�����^1�h�?��cO r�Un��E����Q��1I�UЂ���Dpv#kk�Z�O��>s%��p���!m�¨�K�l
�>V�d.��F���	@g�f'��]Ә���;�*�Y��`�@��O�g7F��������?�4$����鍈@:JuJb3�&���)k����p�
귫�5������rQF���vZ�Ѳ�9A�P?s�bka�_����>�+>���!����i�ՆN�+�dT����X?E�����+��_0����N��@��V  _����j@I�?+P3��y�'"�fҶʏ�不C_S�Y�%�DQ�(C� AtݿgUY��׋��#�*�1�O�t�+��,�'/� ��JQwytWD�a3?���%��y"ذ=Ӱ�(ڍ�i�x�tĺP4d)��9ڦ�U�u��͉u��[B��c�>�'�|>6��l���K��^o�������ċ�Ŋ^�_|	��)��c�	l ��$��x54F��=xm�ײ5؉���J���Mجg�8[���G��̵q�竏�KZ��^B��x��~��{�Є)e�h�I<1qs���?���˒������+OC�c��f���_g�Y*�H�R-��"�Y�����Y�sp��~�蟕t���Y�T��1h��Kbz���o�+x�������+0�LxE�ዊ�}��t��ݝ�|X���H�ĥ?z��lƖ��S������k~���[���ڮ�q���	w���z媞u�"���C?��v<rB�T�~���^���j�f����&�=����)�v���x,�%4hK���3m�OeY�t�P���(K�"
�h��G��Y�)u#d;c����G(�Sz1րϣ�v�	,Pѡ�Dй�a�2<t`t�!#�2ȷ�y��K_�u��'"�P�|e�8�ۖg�h׸\�@dE�|�Tk^�M&������܍�����4H��3O���9󽼀�b�`�S|�EȠQ�fB�VBo◤�۲w�E��&����<(�@.n�U\�S�.��$<�6��D�idJBl�aTJ�ܤ4��w+\o�E� �͌DPQ՛:��C�Kmq�ms�_��P�{.1J�*��ݒ,p�uc��}�l�x����b t���ϙҷi<�eU��߾R�+�[�,�lM� Xj;V��Wg�����%55�~�2kS�e���Y>�=Rs���FT���JZZ�o�(��ވ�+1&��_���w:$Rd�F�H��U������~iII�\��~R�8s=�t�5�2L���N����?�`*�@,��Q��]]���^�~�����v�V�{��o�ե�9H�'Q���uiA\4��(�-u}%��� �  ��>Q2O�� ĉ\��>�
L����;W�M�#u��I6}�>�yǮ��_� �W�2�+�*<)	��L�Ǝ�C�Z�]H��0g��i%	���ܤ��|V��|Z��)�M.�M'�+���H�n�f�01
q�A��ZB��� �� �~���T�U"�+�㒀Z�d��wQ�r��E�rRKީڐ��$`��Ά�Α�Xeq��x��M���Rj9mA�?��6��9��q���y����D�� ��B1L�zIA���Z7�������؆P�[��*��2����Zk�-x�I�6�J#��oKm�1[*�c�	�k-�p�$��V�e|R����4]����a�=�����4�銾� u�R���Ԕڋ�[r޹�$M���O��|�z�@���=��G3]�xrf?�U���K���Mgs�K�r������3V[0j�L��x�PF��;d�~	�}9��k|~#=��BH��)����yvzD���d5=���A��n�t
V��:�����S��D��l�)��
Q>[����� [;6-�� ��~bO�FK�%oD������)m�3����;�"��)'a<���������80�N;"��A�6�i]��w
�~r!4��$�[����Nne!9=��1����K� ���#YY�!�>�`�Ӹ5��`�;�7'Q��"��r���Y�K�V���Ý|����:��7�v�<
����3�e}�,�.[�� {�|�E;u�cƊ�0!fp�Ƶ]��y6>ϗ�E�v��r���#VO��ā��1b��e�wXd�A��kY�)S_�\%�Jw�E�,�j���}�b5~��
��t#U�_��lA��~�p �d�
X�%Ďiw�{��@��뱅+�$6J�BЉJ�$��Lv	2���0� U�J)�"d!�]
�έm����선vz:�n��_����+ȷ�L_:�������K�_ņ7��qH�#O*ǘ^0H�q��s����t:z<TğD�p�ϲݳ�f� �[�*KC���s{��'KW9���;`>�c�M�_����U���q����>Ӛ��\Ѡ̴ޯ����5tP�E`QB�J���\<�+�^e^|�Ze)�� ��^m��� �:�&��,t�3g�'V��R���I�|��ҵ��Py���h�9��N$�Ѷ�ш{�ę	�pioC~��_/��B�VxG��/U�i�C�~_�����y�1��F��#���2�M��'�5|'�P����W�=��3���j.�����ů�Ә�ʰLa�I��]V��I�s���`fJ�*[$3�����cg7�M�����c`v ۳����ɰ�4ZD-���RB턔�.�GL�ask�\�۾)n�_n,�Э���j���U���c�%���΍}��!Ek��I(}�䠀����D/�425��i8 Ӈ�AdDcấ�������j>�����z� @��(u띡@�I����d!�Xء�)�J��]�"u�qE~j�u�6�������v��6��*�3ê;�᰹D87����X6-R�lJ��IG4�� ���̐8�� r�ʌ�zb�]ꚓ����08	�����p�<�۶�6�oϾb�3��ZL�2�鈍����rA��}'+��d��܃ơ�zkr�$o���"Y~!�	W�G�� �Wp�cᕬ��5e0�����M�|D8���&���r��wjǺu�k\� ��,?Ex�N����{�	%���Ӱh�E�ǃ�A�I)�˄�澸#Ss����=�R��`T{����� v31-�UT��0��}��ŭfD���!�u1z�`<(J�~�����[�X��9�p�
��o-�X;1���"Gc���P��p�[��#��k.�$�F>�7U��})~y6���e�8���wd�{2?|��9ri��+F��>�c�*���ХS,R��쏡�aK!R�PP�LH��H%$�3^�s��?|�I��Y������ٗ��m~���)�sr������Q�	D;���㘌(��g����=5����bc�0�Q#����,��nZ���h�����Ǚ���r�N�D9�enD�v_iH�
i�WV*�K�1c^0���D1�ۍ���	��oP$q�'u�n�c���M�)P�B|8jG�	3�h_l�c��N��0d������Eie ���z��"�6�{����D���TEqnU��x������XG䗕ZW��[y`ELfc_D�S���/�Ԓ��� �ρ_Ff����W���\ �+W��Px ݿ7+�Ѭ��F9��.�5,��j%��3�jȭ�l�U�B��v[y�o��+s�������	�_
U��dnY�E�)��귧3�S�Κi��8�n<'$Liwd��&zg�M�mu�
�9�'��G|{Jl=KI"
�O�����)�P�R����7|x/,ͷ6<xJ>��*�c��ͷ�"��s�wnr�-ƒo��D����
�p-5����?�r�~��w��{����CL����H\>��q�����'���xw-�� �e�N���s��d��}��&oJ�:i}Koa4Hg.eF;���#��>[��h����i�r���<��X!N�4:Xw�����~da~[�7p��v'�&�;�G�Zu`�ac�J�!ɡ�+|��'Ĕ������:X��xy�Y�{(���nف��?�/#k��azb<�3�i�VM��,<�x�FI���@�n��L�J�ٚ