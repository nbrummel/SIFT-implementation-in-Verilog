XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R����Od�+��5�k�<у82}��z�GeSH7>��?sEN�
F_�<�]��ԃ�4����@y:s��4O�:mr�Npr~ ��{�3����`pN��$���?��Jxp��B��	�Z����}R�֤��qm��Sa^:�s�6�f=bJ�!(����%k�f���eF������簡�����W�����}�Q�g�o5
&�r:����@z�#JpW� ��c�+t�Yl1e�_�v� R��B���5��&S��~�����q ؂����<�udH��.�Z�+�lGj
��Gm��YrF2J�|��x�f��gę5qx5���	=i�.A@9���Q"iK5�Q�oZXO�i�����Í|�k�
u�^�;U�?�)�Q>�c�&'Rl�qF��d8��q����!盍R�/�Y Zђ��@��."�8��綗�γ�抔���)�W�2�/���gF>��;�{�_�W$�?�cJ�>����2n�'.�S�E��geL6b|�]b<+�ԇ1��(@�� ��icɠ�l���t�k�3��q���)q��qy��T+�נ73�
����,�@;r�����i��Z�7��.�{��a��N��S< �6-z0�`��ZK���u��ߦ��#�D�k��J�oJv�b���O��/\��~��kx��*O曧�V����<	G�a�w���$/��z��(Sm��&�U���E�F)� 6�jha��j�(�+= Z4-�j�7̀���k�XlxVHYEB    fa00    2030Pb�,�m���<m����(�?S��>t(zb���v0������D_�;>�p�޴�+
�G�njְ�}y����j�zE�kRK��Ѱ^b�E���	d�d�_d�L��Ɔ*i��Q��"$Ǎ}�5��Q����=,h���ſh�8�%�"��b��Xi�Z��K����FjB.����ۖōBxj��N�~
�g��ߎ�)�� Q_>�ث;���{��o1"P��d��}�}�7��+���S�]yĤg��لmS�����HXO���R�i��NQÕE����L�� �7&$mvne�9]A� �62��L�%>��?Q2e��9�=�&�oJ(�9�#+N���j��u��_xh��<�k�ΐ,����\l����/~@�}��ǂ����U�o�p=��i�=-�r1��"���VKڒ�̧�c�����p���G�˜#h�c(,ʿ�s���w)�ǮK�)��]jg�w� �f����L�7�:1jn�a[�z��,lfDp{�(�V�&4+���EdL� 8���d���-^���U��.�)��>�����g�K���$�"h���&<4�ٍ��7�VuM*�6���D���E��9iw�O�w%���n���KkP����l��Zr�|�?px����S��\�C:�t�2��R�s[zvD��{>���Xܸ1��)^��i�9�y�~�65<��Ҕ[��(	�'ؑW����Ehp�ɀ�.6��m�cR�t=�����6L�`,�8�sb�k?������'��H�i~IP�=���V��f�́����7�Q�� ��ॷvQ��gA�軶��%+�RL�B�l��|8B}��U=��'�o���j��v�">I(���@1�	sZ�E�x [��i�
bR~t��~�Ø^yj��fv�v�_O0 m�bb�g�VaVio�_D.�MT!�#����������V�t�q���<��dV�x�g���*h6;婨H=��-]�͡�55��(l��.��P�z��pp&+�tZ�.���Xr�K,�8��0����,���A�Ԉs˭�D]��N	�PU'���D���J�k�P�S�tDrZ@يб�9n}6���؅/k��c�S�<P��C7#h	��.��F��8�������X��N�U�L���Ig�{(_e�s�:B�k����!r��I�nQ�u���V숌�.��N��^I�H�OK"�i���e+��$	H���Jqza�t|]=(%��Q�j�pw5�vab�;�9>�g���RX6
�x��&\C��2w\=M�n��'�;�VfC�W�ʣ�ʢ�(��z��Ve5��5�-��mK �6�Yc��ч��=��fD�^�a�d��gUd�Ku�I0��8�����zd�g���ö�\�%(�4r��v�[88q�����8ʱks�T*��Tסּ����������&�~j�)u�{��<.{ў��^3�@����T� ���I���) ��(��ؙ�6vܛ��#=����v���c?��u����4�qzc'���OJ2�t��*+X������6��]F�7�1�	�S�f����Z���IO��rt�i�e�=\�)��K $�3�^��Au�Y(0L��P���ʶ1wCB���#�s�  �6��O[�h\�!+7�� �#p`����Z�*Hn5�?���A���B�.b�����
X"e�eë`P��`����7>6�n�*��8�2�l���]�Dgxr](4F��p:��ϕmԄN\k�
�M:O�i���_i�sv*������M#��
I�ȁ���m��/�g��zU6>��������@D`�#&�n�
|`p�{�W��,��a��ih:�6���[��QZ�|� ��`Ġ#���|6��x1N)�;��s����t������M�ۣϺX��'V��Ms�z�>ڏo��n?s�	#YA�w�A��[(n
�	��Q�������*�+�x�)
U��`��r�H�޾ťolA�ې�߱�N��!r%�n�]����8�:�}kɃa�6�|�K_:x5�߂��4���kf��mA�is��q)m���	풧�$u<xF���^����<�)M��vƨ�j���j�q���^5͇V���h#�6�;�| f1�}��5t��]$D����?��<�_���j)(Kr2C�,�[����Y��zK^Y!��ن*�|��[Σ�8�X}�Kk��[ϙ���� ��h�aH%�C�����!.�w+϶�.�OkKc5w��N�rX��Ɔf��O$ITS%u�~,&�b�W:ks�mD� mׅ��ب���r��������4nzm���	�h� ��G��,��A�[��^B��)��h��cDĵ���Co�`�� Qaȴ�(�l�N���\87r����0�x5_�1Y��LS<��q���]���{�Vb���07'ƈ�=�2:"��	7@T�1�)(-��'��}��z�L�_�|]�ۧ��� �߃�~"�|y�c~ۀ�Jn�#��}�k	�@��*�`M[ �)@i�*�/QN�C�z:�,�u��&S�˴L�q��@��t���-���U�ͭ
wv/޸,�����j2��r����D�T&0�0�"��t�<�鴑4�@a�B%�Z-�~��K��!9�����?�c:-��LV�js~#N �<۹>EW�vC&M�}Y}�$�,P�_l�uԵ%U[��І/�w6���ƕ�H�YU���_�_YH���v�w��_9�dx��G^pGze�G5�m�oD�Z"��z�?3r-��Q�lq�S��#v�K��"fKQ|�VoNT4!z� �Y#݁z�>�p����vψN��U�nh��,�<���R_zLd��w�����n��]p'K�7��E���-��(i~ʟ��Zy�b:�G��{�U�eF+0�)�n�����)�1�*snR�co.�+��C�c"$bl0l����+j:���o�+O	w<�/��+�1_L{��hQ�l�f��5���V�Rs~�&q;ؤ�M����h��m�x,/�صۧ�A�vxQ-	���"��r��&�ۿ�P�� 7(n7J��Z?[��D��U��Tޙ����Y~�u�L��U�Kߗ�چԘ�hS(Of˳�
���C��Ƕ?KM�F\� ��x�\�+�Y�'y�]�#���:���p�Hx��2D��p�P"A����!t��Yn�q_�)�f7h]����F:��h���0�,�I�|��P�� =^1��G����K|6SNa���`!���e64����C�Bn@%bh;��& ��#4,�"�eP*R�L+�� �7�}2�qn�JF�ֲ~��6*�����X�ũJ�
 Iܘ8(�L��!	t�"�и��I?r��)7j��}�M�d
���%IO�%�<����ը�В���TD&��!&��\f9����3�es�o2RC��Sԍ�g�D��$������,��I��KnV�ԱOfUB�Ϯ����Ɲ��xjˁ����܁���U�箑�G�L�����XH,ӸF��/J����5�׏��j��	���c�" �p�l�nԄ�󦝩���'!�-z�}��ԩ�f��M���;�>ˁ�:r�7H� �O��xV.�7>�K���_���`�b�E�-�|w��"�_���.\~Gq�HC6���9L��}ص���Av��d"��Z ��������3Y��|�rJ�?�aL��Ʒ�Z���N���UP�=��R�� 8xrx{�� �����9ȿZ����fE�w�^4n\��j;�	9n�>���n��8%��!k�_L��d���S���<�˗'�1��v��9��7A7j��N4�`��	Q�Pή�Ӧ�~?�c�\;I�h�HC����:79�������@�Z���N� �l'd�K�lKo;�GFF2=7�~� ��!܅@��bL{�4Wƃ	���*��w0��]����D7��J�s_4P��K���a3��΂�z��9g`�1�1�d�3cn�B<
�|]��5��	�Y'CN�Ol��'.����1�����23�:��i[K���Q��R�0�ڗ~F��F]3'd��U[^�}�|8���R�^e�T2z/�qp��-�+�%"	����aDUB��Q��9�f`ڙ�&��d��wWίi��_UD�$��e[���C���Ct��zJ܎�R�[�֐��Bt��K�c��ɧ���%��B��E���L�����}���؏0c���2��w'(ߞ�� <(��楂���j�����_[�l�������J;�]J;�G�rxC�|�r?��tp��i��D[��)EFE�*f��!v�N3��A��T��>F['R�n �>D.>��)�ݺ �L�{�w�/gos@��8����xQ���.���9Ą~"�Q�������`�/Zx* v~������=m���7N�5�e�`��N#���U� �zH��mZ��Т� ��(X��$]���L@��,e�v�T6=ÓS"���iPy�����e:
Dl�a�c�^x��0S�a�O��ώ��ٔ;2!�o�sH?0�6�>Q �vY��`���������;�2��}�܂eS��H�f�}�8TH����T6,c��!��f�d�S #Rgs\�O��t=���"�E�8g@w%AR����B�]�O�E�њ�B���|�=e�z�#g�VF�����N�����W�l��X�y��� �G��-��+�,J}���N��;����p-�E���k�(�_	0�=���X��8n4�^g�6���sh'��iu7�
���?�1'q�qo���ֹن�l�ť}s��ڄ&j�RK�1S%j��R�����g�X;t�rK�_�{��~�:�IO�˚�	M�"fBʯ�9Dxy�J8J��T�2�3��[�5��r&v`�x�{����^�_��{�f3�X��oh�L�AZ�9�"�&c۟|^�	w����`��eM�*Le����Q�;����ID+�0�v�����y>�+��$/6�/tEJpS�ݮ��Nʷ��de�AE,�����.]sh)U�h�b���	�L|ft��5�xl�z��`��m8&q$><r�$*��I1u��њm�n�2��5��:�?�}��R�y���E�=���k�U�L�\� �*��^X�!�&�����y�L�\^$�а��;�������o�}f�_G[b�V@欴���%�xɨ⋹�4�<85H����Ӵ�ku�v�YPP��Yh;L��>Y���%:j�uJ�MU��	�Sc8���ś�EA��6���ʙ ����)�1a��B{�|7��(,���G';c8�+	�>z$�;��a'@3�ƚ(SSCY�E����:)ة~�F��o%�]���җ�Sh���nD�:�V���aM=��~��f��49�g8����bRo�a��^fp^�K'�m���T�%\�2��� ໃc>LD�z�!�ꐖ��?����i�kJ���w�d� ���\Ox�
�+����K�(W�I��\��׳���;����f}�n� Z�J��i������X���h�3A�*�[���;{:�Z���R�RXC ����-9��آ��A��p@)b�;6��*V��TĶ}����έ욦ӧ_AT���P�b}���HB�����z<N9����	^6N�l*���eRbj�2DR0�ǽ a�YWuͼ�-5,��U�]-����h��a�ϼ�QsP��R�LeRݟ�E
��F�Kiy�~�[�d����|��(�1�'�H�`B�r��x��8���b^2"`R��Z��w��{mӀ��?J ��}���$+b�D�B����\�u0���a�xԢ+g4.�U(�e�ѿ�B�=�{Pkڏ�d�M�l��,�$�-�i�,��*2��ۏ�ץ��C�C�`7�+�"ӕAs��ձ�g��~:ղ/V��J�|�`��6��^��.�?1�s��9'��|�L��#ϩ��Y�U`��z�n?��&�Ì��<FH���IOϦ���5>(�8��gv��N@�˹���^Ƹd7BV�i��A�9+��v�R�ʝ�՛��\<�n�h�vf�~-
���D���Hie���>A���`e�K]%��������]�e�.�S�j�3����fNm5�TN9�8�x��]�\m�Q����[9 TeW�8P�ۜ�1���S}8�b�ݷk�$��r�O���8,4��L��� �q�_��7MX;>�=;�+�����3���K�\�K�pQ]�k��:�!+��*,F�ܐ���,�Ȍ����P�9��z���y&U6��P��2���z� ����v�Y�y��d��xl��!އ��XIR�D��%�������c��.d�6�=���h�&�2B�oZ��\:�bI|d(O�U��42/��^��D����:
�7hɦ�N�a&���]�1�F�J_h$��L��6Oދ:�?U��;� ���^M$w�a�A�,ŉ�U|*�BZ7�i�İ5�r���$R\s��@�H�f*���F�W�8h�ly���ܟB27z�=���->k���y�S�)�-I'r�j���/���}����B�~՟��{�ƲIg�w�y�JB�KTq���Y����-���0��́ڱB�aM���1���ۖ��ͺ�j|�&9������L����bt�g�?�y?a^!��j1����M}���ت���D�Q�L��$Up�Il-����ɳݦT��(*�<��<\�[w��H�+?K����"U.�]���6��R� \WZ��$�c暪�i��	��ܟY5��}_|a�H�ٳ����c�@�*1��K��p�>�����W���d�;E�ڡ�V�K��&�١��ʿ�}�?-��n�s/���eP�k\�ӟ�'����x�3��B&�u������d|Q�@�A�)9�Z�iUr���s� ��,����w�j*����Ro�#�'�Nd���4]ez8�h����uJ%d�n������mO7�^��)�b/S2�sy��{YZ��8p����O�9�Wu5�����P�7��9E���$��5E�It��%|\ݧ'	���И���K��k"4z''cF^��B�f-�U4{q�K]� t[E��@]̍�TY������m`���<�{�hVa�`��l������|CH�B�S!�v�@᜝�{�9#h� �;���e�{���(���O�\U���^����r�T���OKʤ!U���Wii��ɋ���ѓ�����N��􉍪t��ӻ��L9�f�l�48@㮕Vr��v����`@s�.�WNRE��A��%[��S���:?�7�i���MH[�CR� ��D�L�@��#-]�y�5�a7[ߪ=�&���q`��a��ʞ��0�Q������2A�=L��cwp�(@�<^k�P,�k6o^
|�4A�~�yQ�`����0�8��J*�s ;���]�N�_�ܖi�翥��~�RJmUt�ܫ�1,�5�����Cu�pU�yz�[�M���cD�3����v����LFV�{���z은�B8�V��kw�X��?�ؘ5�;�����U9Kx�5t�f���mY���m��A�̖	v�d�k&ar�Np�\�����O��L�R'j	E�ztҥ�dag�u��b��Y��+a�:3 ��!�1����E�a�QE�m�i�C��":���
��� �%Ԩh[��� ���3��W��p�3���:ٙZF��!�G�%cȞ L�uՕ-�C�y�
�<	ϰ<�z�1u�631ʊ��?��/$p��^'쇾��,A�&/�pA� ���[�C���"�:mN���*���"�M饺7�9�J��L�?�iqQ�e��!.�J<���L�*Ë�h�A��>�}��s4��%���}&��3����,S}����\N�B� �%,,-E#ס8���-bs�B���Z+��`�"lq�_h�S.���(���>6��g��	���z��f>Yc[��VU��	zx)X���w�,Y}������c�cZ��rP���pr;���ʼƻ��H���>f���3�%�;{,�m�!�HPQ�
�Z��溦=�=�A�"��}rAz ��ڋ1W#IM,9MkҜ+� ��ϤK�?uXlxVHYEB    9620     d70���7���4���؇[G,������P���4����H�+��XB�� �[�?pN��d�K/L9�N��Y:Y�"b-B�2�?HMH����u�:� in�Ϊ�N·�%8H�2�M�xA�n��X;��ai�&�цQ6��G K�ȝ��0.�3�(d2�6�j��!���~�P�qA-@-�B����a�*s�h�9W�M2`�jA)� �9���YT~T_�
՝���`�	K�Pߖ�QYELu�|9נ+)�E��u� �����^T� ���ZiJ�Ÿ��������=1 �;37Mv�2���vw���4*"�Sf�Y+.��fi��"/z��5�ޞNԱ^��}~)���Uj0�!�$�z��\�\W� ���=�{p_�;��f��F!�\G� ��$�t��j�4>,<�{��v������?����[#��X�B����t=�*;%(sB��w�8<�d8�t���u�&��c(��{���;]���e@���B�M��T�1X~4��PC��-f�9��V����L�L����F@qL)~ʖ���1���R|'��Ӝ>0�%l�N�%��,�Q����%S��[Đٲ��T�6�!�+�!lq�����ٷ��-���!/��nֶ#�t��BU0J&L�^�|do�'�,�[|�1�V=�����"L��7VS�(�ug�  WBJR9�@�Z��/�d� Q�}[������}A�]n���g9����n�Y:�ݵ!�>�p9�yv3�T*,qmSk�+.��2�}�J՘�g�������д�L�
4H�#�6��c�x,��lZ��IC,�FO[�%A�P
FŲp�Lյ!�~�W�U���@\n�m
 r��U���C�p`�{7����UnFH�e�e������PA�/��O�|���T�ю�u�d�+iF�z��ϫ�����5���̘�Z�+�0��D|�:&2��0i�*sh,0��������H/Gy&c;��"=��V�5X�c��=�f¤�K(m�!8�@{�TO8�������{=&/���I������� i��g2-���`���O�ӌ�SWw�ϻ����WH�3����8D�k��n��x�%Q}cy�
��q������#"��k��*���(���P%Z^lhu5W��J �������v��Q�-���� ��R���qk�K��T*�ļ��^�ӗ�P7��kZ���$�{���ڎ���T��ڗz_�(��5_�f	3�|�<!�u/�cT�N6@=�0��#B�2 ���:
N�y|����wS[a�^�[�auY�g��֗��?�*�8ա�<�{m4��<)��h [��6[��Ĳ���W?�:Ib����Z�����!Q�P�F�Ж�z<�$ܛ��;�@[� \��m�d��2軱-����Yݶw�2���I�����&V0�U���,������˥ĺ��%o�Z��!E�������Њ2F�X���tP�!�ip@�e��	��@M�@3��5����S�IPOM���m�=�LMd��5�C	��,� Ւ�����!B��\�L���d��G��э5p��_�w�N}:��ӛ���� �=���^So���J������%��{��1��Y���]�9�TL��<��A��{Tϫ�Ovu�O(S�a�����i��n�����jz?��_n|_4<�K`z�֪4w~4�t�p� r>�d`�qv��M���z��枸n$��T��[ �J<.�pF�3T��X��k��K�{�� e�]��ׄG4�aW[�V;��z(�nu��,�.�Z��)�WK����L�KO9�K�x�X��sg���r�s�e�c�} ���v��)V�+�;�$��W�7z�x8�ŷ5������Q�J`���b��\�L���5�e����^����o���Kܩ���]�v������G�M�`���͠�m`E�ڪh�ճ5�۔���p���>�A؇?"�y��.�T���;m��E:^���E�hʇ�9M�b�&RF=iM[��p'YMw)R+r]M�e4�*5���qS
6t�y�����h����>#���n+�H1\
�=���������g�Ѱ��p���Nf�KG�3���k\̗��t"o�SL���D{Y?���Aw |nO��.�ߜ���Z����Uҹt�[�����@�Bn^��u�7�kI�Y��"3���vpF�m:������{�����#B�g5c���K�V-��~d1�[;	��Z�:��~f\�c9���f��M�z�8�
��Z�[G�����~�R�uBb<�U�'�F>�F<�~��%��(�p1���u�C!T��_��d[m 3��04����/��@�m�N���A\Z4��w��[�4<!�݇���T���eŏP�4k�]gs�g�l\�f�)Y���(2�`uM+���/��π�#�9Ue(*4�ѝ�sI"�ӌU>���o�i��*�粼���{J�����d4��/�e>7�E#~��(�*���4���^5���ۃ@��J$�����d�+�H��'Ą�*o��	J0��̛
c,��9�>��f��PE"�1RN����G��,�!�Jo���y��5�9X�?\�26Tf~�2�f�@��*��ʏ�����u��f���?�،"�,�e��8t�S43q���}�<��H����'��7G����g���H2q6��ӭ����&��xP"Z	������wo�����
$�1����!�����E�P��:��j�")�3�0�s	�J|k��<����܏:�`�&��&�2�/썸4י�N����ѻ���Z�f��=�� R�*�P��:P����~�(q�R�c��CWS/��ͷq��.n�_�'�@!wO���5�-�%e�`� N���H���L��*�R5�E�Z�.8����\Ȫ"����,��2�ʍf�c�t:�+�#.3u�׹����Ǚȓ/�}����^��9~Hq
-�i�����V���<>���>Ī�������m.7]�Qm�̭��:LD-.��f�C��4�j B�|���hT�f�w���Í8xyJd_C�I�tՑ�I�3��Y�9P�Ѝ��[��LQ)lN�����6��콧W�PծJ���v-5��F>vk([�Z��rC09�@*�v2�Yh^��M�B�� ��)�I��Z1K�k�>6I�a�� (��ڧ�G5�In!MC�-,���#m%4�)Q�s�z3́�p��1�D�U�BQ_[���o�����^d<QN�B }���a���U>��ͻ���a�� Mx�,*�^W2�/{���� ���y=X��&�M�R���Pl�Ig���pJ����,kDT�-�Q���