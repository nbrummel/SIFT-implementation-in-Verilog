XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|�?5�ݑ�F'b���i!f�on(�ߥC�����a���R���;$�x)�Yƚ`�����W�j%\8p-GƳ�#������ 0ݴT2��P�k��.���V�S����	�W��y<_��Sd���E�dkO��P��]���=%���_�����ĕ2���5�Na-�r��F��H^��	�(��^�8=ӭ^�io�H�쳤�\�a���<@�{	�l۳7��.�}�E�Pf�;?�;%����{���DTo���������E��y �G����'�:�x%^HH���w	g~+n��|<Ɣ��l;�i��y���a3�I3U��O�j���	����d"�u��dk��vR7����i;��yF#����(�,tO�k��Z�V�ܯ����������&���-�>�;�G�v�$[36��T�1��Š��u<aY�����%�;sA��4v���p�d�}����>�S��f��{��xr*5F.�p���A�܏�Y�?	zCmP`Q�g���;v��z�U�Î�W��W���^�4��I� (��z1%��~�1���й`���k)AL�u4�,�s��ރ��7x���|��;��
��s����\r{q���<���w���1KFaw0�.wn�(����9(�����
OH���9B�T�����~�|�jZ�'ŧ����x�Q����I&�Ѐƙ���K����eԙm�����~���[c'��Z�<u7��P"l.��*V�ڻU��|:��Z��}��(6\b'XlxVHYEB    1192     750�#��(%�z�$,�!ÇY����'�������[,j6G*��G�(��s踗��qbĮp���j��x�~���my�&y^akNz�-k���<~~��f�]�q�)>���pJlF���ˏ���^w~*���� ���`M3�`�\Ly��F�+i�,;T����!mɣEa��J�������ͥ{]�Ǫ���E�t$����;;�d[F���zK�7��\p��_��L�p�������)�S��1I6PTjC;��S��-� p8�vG��<6?�������P<jڷ��fX�фM��!	�����f�]�#���OazwPn��Z�KV��q��fB�#�5�5))5|�uli֍��_���W�Z��µ�Ul� ~���g|��Z���y�p��bg����b%��޽��"�a��y?;td+�.6���=B0�����T�l��;D��Y2��=g�Nfњ9��׉h�B?-V������ê���n�/�q�wHI*�Dv���y[2�?���#4�ya!��(�嫼}���D0�]f`��:[W@Y�,��S�C���� �m(׏�٘M�h63UE�vYm��.�b�������Bq���uV�=3�
�"�#���o��w��(c�^0�d��KDy��;¹�L91����#��+�3qU���k.8^�,��:�{��V�o��j�tQ	������xH�u
e��ۚ��y�Y�3�u�݌U�tQ<V��oK̏e��".`+v�Z��g����9l/P�'��dԙ����Y��Jj�P��@jf����c,���*�A�TU��s���mT�ڦ������A��a�����K���~�zĊ|�A5��H=�� �v'�.O<�x4A����Q#�>A�t�	�>��iL�|o�|J:Vgp�j���g�Y崟��>�7�0i���/��%�����`	�t�3����y)�#��4�D�����+K�����lb!���LK��j3<gR����lܘ���b�E\��U�Vԇ?������RC�^7��$|��^и7^Y�1T�j`���<��
����r*�oŕ��n��f

�p�BTM���\�J�lT�R�����yk�,l��I�l4������ 6��4oOY� ��ޕ��Vj8�I�LF`�D��f�"���$��=N�>l˽�{��>���� }nպ�ŭ�o}�>M`��}����М��mg���]��(/�R���9�H�0S��̴��ν��l��[�nt�3��M���*uSس+����Jik�e���u��.�kQ�t
sn��O��n���P~&�6v,��[6sm�3r��6��ZB�z�]��]4_�þ��''��;7�������r3������1�'˲��T�f�(Y�c��,��Q��rf��#��o���T)~S�}�.=DVp���M�F�%�0������Ax�H���[\56e��rjH���bwM�dM�[���
$������}2�O{/�^b:�P�DM�P5A�Z�qC���o�e���%7ZaX��G&q?P�E/:kL��M�Ԥb)'��[i����r��o�5:^�ց�a������ƭ�<&�\�G{�:}��sZ{�k�̗�qT�ῌ3��0 �F䄝�G3YOSu�>A��ic��IQW��ބ#���C.���|�ˆ����&=��g�RY{�F����s��"����X�z�=#��p�q��Ȟ!�dSY��C|�^|�i2j1v}�'�Pr'˒\��(:�P7�N���1S]BvY���j�}�>�_��Fe\��WSѠ�c:�����ѵioW�~hq���#�1a�}���jg�SvN-�L0