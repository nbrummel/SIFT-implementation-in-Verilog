XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����c��&����sy�G��.������_�$�C��O�v�]�Q2b��;�Y	 �Ԩ*���ȞX�=O��k@'Sn-��	���'��?�7��K��6�[�����H�+tJ����	ՃU=@�H[v��,/A�P��;@r�%^�,�z��!��xƪiG���
L�l����g�7:��Wwb� a���6�e좯9wv�.о$d�32993}b�mv�� %�Xh�aN���`斛��)��A"VTw,���Y�{󠂏��O�S�Dhr�{m�*	R�Z�>�c���|�	�i��A0����~)������#�k��*��M.G�����V��B3��t���G��+�1����Be8�&������\�8��6���g�t���L=�f�z=�����_����?V����"���<����w<E��oZ���ze�"n��_%{n��N����i����5-�n�1Ŭ������9^�\~B{ئ�n�Ț�S�yŋ���76Ţ�U�x��̣���K�Cj�����O�Y[�*kN�&�ju:��ʢ~��-����~����+B~I�9��"&s
�i����:�|�'�״	�n��>3��I���x�ET�-a� �ۈP���fU�<^��RK�M*s6�
�4W����#~򓬿[���?���r6�Q�(���v]b/ۭ��QuZ�Z^�"�pf{C@MF�7ٚg��b�C���F�y��0���B�O�B�@tw�j�Ib��<�XlxVHYEB    2cfc     c80�݌+�j������Q�{$	}��&ʟ�bGZ����V$��ذ)}c�Ǫ�?G��誠�载YX56Z;���MհTmb�_'��5�K��q���([/g��ک�,��@����'�zB�$���� ՚r4��N>�!���.j��%+Fj�]	�l��ۃ��c=5^����[����{E��1��va�鶯8k��h<�A�q�lc��(Q�B`�m�u��3��р"����G�γP��n�Mcqu�%"E�n��'>j��i�4��bj�]���׹�z�ߥ���S�v�8�{�)�[2(
�����U����#����dIgI�"��'H>Wv�����zd�EԆ��PW���⏒�MSk�|C��usR�F`m.!�W�B��#:W	>��}�#3,��o:ѓX�M�:]�jP��0ˌ�(� �K��b��9>����K���g� @����_�j�h5>�zI.�(m��Yr���S���T%�gkҀ+��3��]tB��H�Vlɒ�P>��vW���*\ǌEQ�/T��^)u~^P�?�@��+���[�P����:Υ�+��������@�����B���P�'Dk����g
-�t�DyG^<�	����JP-�"U��x�g����[}��4+|D���	Iqu��?�×����s��|�=@�'�A�7�>�l�(;�f'��s������k�E��vfo���|U(f~��-0�-�l�F���"Y�K���4.K��S#[
D�������IbY9����{�CXp5���>v�o�o*Ve���&]N���[t�U�C����A����i0Ga3E����ޱW[q$�|f(>���?����:�cL�΁���u���Ӌ�4�f�aK�A�yx:�7�N�۩��zms~��!k���=t!�s���4L��G�E��I\)xd�8鼿ݿ���u�[��gt�Q��	��R=����~K?U��*�3����w]k��_�z'>4;4��y!�3��k19B�{��b�9M�~�:0�u
 ;�vؕ-p���VW��I��/~�I�]��_j����o��D��ϑ��M�&�1���;�(Jҏ������7�V:)�Fk�3sf�s#Eq�̋���{[�Q���:�E�=�5��z54�-`�����m��%��+��#�=��t�=ǒO'�!�-1�����٠ɜ ρ��ڈ펝O+^�dZ]��B�˶ED��<�j���B��g�KR<���^��p}����� ��CC�4	��I~?����6��>S¼��y5i���H9:����*�t�]H��ZK�S	��Iǩ&����[{5��q�������>R���gME�|�H���J�J�&��J�F5Q5뇞l ��0��s���Ux[=$#�
�ݔⶶ&�[9U�G�RM�jAF�qߊ�7���T7����d$���o��r\����(`��~]�?������o=��{9)'�>ԛ���vx�OTp%v�q)W�6�����S����,�4H�SM�k�=�_uu1�?k �m����P� O~�F	{�r{��<R�(����Iu�e:�o��mm���+(@v	�)�[�y\��0��? ��dф�k�?�(J�+���_֏8�М{�jO3��|����������P"��6�&�%"d��)��q6���8����$&��V�c�N0ew�4oS(ߺ&������l�(8(#��3]�~�x;�4�)�Z46G�r&�>�9�l��/}�q-�!V���JN��uï�-���U�ZK�Br~��3<޲md��'|^!$3hd��-OJ�tOs�+v���n��ʋO`�����;>%��6u�[Wx��V#�S�4�p�bD'E�115\p:�QImBG9���*a���>g-�k�-`�Ƹ�2���P^�d���Vp���++�wU�(�Z�}ϒ�:�\t^�`L7:�ӷV��\���,B�G֠��B.X3#�^s��Z�E��+����	o ��pH?wTÇ*�eE1_%�lUe�C��H� �"�d+̙�� X]t$��)$��J{��a�ꄀ��F;ԍ��Jd:EC8�^��x��
��c��D`Hs�9�ȩ&V@��A4�iQ������٠�-�*�H��ݘa�������ru��)M���'k�jyh��%(-�@���|赁�[rOQh�;��tⱅ m �s}SQ�U��*�
�[.�2��w��{l^�OM����%��`��%9��r4�4����-Գ�Z!D��70%���ߓ��
К�� m�e�Q�8�����ˤx�-#|��c�*J�����3�M��f�tG5�z]��3�e?t���#��a�*��&8�\l�P0���vC����9��{@9?�0�s�X!m3��՚�bWYPe�Kpq��f��Kb��Bw�����Gm�M�.{�)�׍sI7�ӢU%�d�c1H���9����u�<"�W5��]���U6�
��2P�T0�R��蝷>����u�nN��o�����'kij����ŋ�Cv��+�P����♩1�t�A��wr�cTL_=�R^l� ����u:3�ꈙ�F���!�>�+�Av5Z�S�Pm����7	�"1�:�ű�͢�ލ�پ&-��,j�)��e�>#�Bb�^E��8^�oN[Z�֦�����״��U�*�����
�ˎ��{�i`Dn]����
(CY�e>;�?9'gP ������ )\6x�����W��i�3�Q�ŝ��U�D�?>���)2@��L����i"T�M�v&	 ,m}�*���7J��uuۇHM���ӿm��K�Eر0�Qs�j�E
j��8��R�w.���I�L��4P��v:И���)�h�ʬ�=�).}��Q���{����U����K�(������	� ��^a7|͋͞	ɗ�K�o�D挟�������a�7*]�����3�>����<Ae�@�a}� ��E��°�����������ͩ�'P��b��YW����_Ç�/��� ������WV�1���7�֊[02�8���c�W�C H:�]�2���M#��i5����>�i����(��#f2�?/L-�fv�i�b��`�v�zNY
Kg����\錄����"��|��C�/7*YJ��զ��91�