XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���I���Ә�z�#*�[eD�y��9=�tk�=�)��y8\�հ��O�!��̀�X�`�{;e6��Vk�y��j��V���҇�~�k�k�9C[���x�१���U�i��P��ݠ�ʉ�����X�3篯�]q�J���9n�~�ΊWu���L+�@h�g5|g��;@mz9	R��u�TҊw��(�������_���j}.u���aLy!����%q��7��o�����9�-d�XP�sd��LYƯ���ڴ��7�#��� w�.<���+��6q|<�iu�?�s�@������_�&Ao���ӽWxr����@7�����W��U�r	��o�����/��Z�:��n��� 0�'�nCA1��p^!�jHcl�`bs>� �(�m���*�[��-��ǡs�����H��B�`M��ءb��\�k���P�$��T�����cC3�G�]�o�nT��A�����6Ů���Qn6��ge%�l`��"�͂�o����ƿ9WdE*f���B�&��K7��:��v�Ź�[T!����J� ���.�x��vZƊ�ƗCc�(Վ"0��N�ˋ���yYTj���2$}{=�	�gs(+p0�t�m���T�o��HSwr8 T�J?fە��=J2����Ceh�B���x�O�,[r[�Y6o��"	جv�v�/����8��#��5���F�� ђQ�~QA K�[��{�VM�)��]�ts����c;,a�N��XlxVHYEB    125b     750��+�+s���х��q�sY$�J�I�~�y�ڃ�4�KdN[R�-��ژ�>�}{���X=��Î�r���PzZ@4�4��fCt�1���p+�o�l�!�żpJ԰�9�c�߾{].�c �o���%6����'��t���Hp��Ai4��A����߉5�i����$�5J����6=p�t�9#3A&��8�5ٍ��*V����/C�� ?�MQ�<d�*.RTD��դ�7���[�&��a�#ih��(v���*"�I�<���ʯ�t��.4��
?�@S~@�����it��C��1��9��{/�H^�Elن�Ѩ��}o}>���wH,��騑t�(�KDv�~ćB��6�rQ�8ӵ�	�U��ι�L?Bu���o%,����oq��KHZz*��Ŀ[��2b�@�_�C�I�у5�	$���ܤh���Ϡ�P�d/l��3���'�r���q*/% �d9v�%��*G� Ul#�\yK>~�A8�	�$��gvL���հ�s�{P3�uۍ��t2�q�=;� T��[�]�Mok@
��ه�JG���1�(�C�4<ڕ�k[%~��k� d�G�X����#�C�ڢ޾�q_�`��$��<xmĄȯӺ�hZ'9e3�nV�1ϯm�k4k�(�?F��xD�k����p#<f8D��F;�ŗ$�9ܮ&��1���qZg*�U���p�9��ꚥ婢��W[Y�/�}@R��1k��*�o^@��
��2�:!��@B-:�n��F7R�@�(Rg4oW��q5�vV�K�p8�x\�*c�<�Oos9�L}�Թg��\�_��!a�ڟX�G��� �
M��f�=9�$��^	�����(�D�K�l�+;?v�r��^��B�ujL_�I'��⑪��
���^4�`\�� �Xu�}*�K�	ع�ʱ:WK���YN�^�,,��)9{{]"2R�>��=� "�p/���;�����Q;,F+��N���i�s���%u��|�u�M/wX 6���,ػU'Hf~��<��o#b�Y�F	�o[��lq]�@q������K}�p*�^/�쫭�(:�ԂS�UYd�g���!\_�`�{^J�`�,;�f����P��g��t��Dِ�y��I���o��"L��#m��f�7b���WG
� �Z/)��B��ob,�*S��U�����>���r�9	�7BI��VF�w[W��ash6ߛLf���@3�3"���Q��������a��(u{��Zɜ�b���eT�b�i��!��G��b�2�MU?%w%��R]r"�5�(at1����@�L`��l%�ؓ�� �(ţ͐y~_u�� Z{6t��%v�g1��kHa�C�:e��������W�|l�(%QaIz�������S�����6g���{܄yB�̆�<k���غ�g{"w�,��!0J�H$�?x����k���EX�*8z)�9�2��F�W�.91��<�2="}7*��\l5���
 /Q��nU��j���/6�b� )�[R�u��}6n��s��i�5>�D������%�6wwRv<�2��1L���&�����b��e�&�����y�9\#PZڱ���2\�|GVC�E_[�����h��b���+�1N�=�W�@�`����4 �y��vw�	m��Y��5�!��*`6#�cR�?�~�gA%�c�R��b1�!�\=�c���B���d]����S��D{��6߾R��(�F��2 \��b���"r�5�q-�@x���2�����:3�c�N��S�$kd�t�f&�^�{�T��q���JP�k��S���\��w y"Jx�?��H�j���a��