XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���I�&p�v���`��y
7f㳻�Xӳw�W�o47�l�V�����EWb�d4s��d��E���W<�8KX,���P
1p�O��
j�VV���s�͌�R<�C�ZPZUgn���=%·!�,��f*C�x�&s��蠷�o� 	~�μig)<���2�-KS�K���]���nD+[m���گv�?��.�7��}b�)G�{z	:�<	�AX���rTA��oc�㪷`�1*�B�3x`�_�`3�w�1��I#D�$i]sݿ�j2KG��)�tۑ1!KT<zf���7��*Ս=���ܾ��EcT���_����j��"��]��4��.��3EK�[՚��}�њ9�ԩ^fO��~tY=^Q�yJc�e���r�R5[��o�S�=�Ԯi��8��l�Lq%��6	 ��V�]
�焆c����o�~Z�����_`��!��֔-o��h.��[�$gU�|\�){�b� �;�댝�"�nq9�-u�_���U�%`�ȇdƟ�R�]���4�?��v�aC�y�O�z�/�V�7�2�:�Xӗ�Cd����r	Y��J:���Q5I�s�mi&"�/̂di������˰��}N���-� K�dfz�fo��`�mz�7�s̄��❺��v�Zv�|�Cj�Z�ȉ�!�ē�Zs7?���`��Ϊ}��Z�:��e;�Y��D����� �n�(@�'��v�@~{v��!��j �C�7T���ޱ�X)2v�y����|���<�B�$�`��Ƀ%�	XlxVHYEB    838b    1770����%�^��rGt�,�~�%6�N�1X�s��w���Oq��9��l�c�m��>�����(�%��5�?���Bh__7�3b���I�ߧ���hq����FA ����*W��m�B3îs�7��_}K���e��"dt:���J��%\��''�o%�"����&Ӽ�e��)�I�:c���@ADX�y���֟+U{U����B��^zzR^�W�-���FN���9z�g7H=��}C �q��1�_�h㬕���&j8��<[��BZO�Q�G��֊ė@%�4-C�89��dJ+i��<���7�	,�D/����pm%W�_�1���~�X�T��Ҋy�`�ȅ�W�5< ���i\�-�fM~�/�����t�Bl� ̴���5����s�GܸFtS���p�.:Z@c��-�$
K.v��|��ԗ��Q��yPXc�l�1 {kT&	�"���4�Y6a� �ۆ?��_�{��P\��'����U����� �VT��u�b��+���2a���`��R���O@3^||.�����)����:��碥I�_������ _�5�TU2��u��}�
~�<��̥b�o��K��F���4�d	�gT뉬����XU?�^P�;�s1�<�pZ�E������Ҏs�W\�4RT/�lP�0נ����]{�J��]��!��O��3Q�֜�&e>St��~�%��]M1H���q0ݯk��<��0���>�	�K�+_o]G_���e��X�3�'�ɿ.l1�	���tѯ�X�4vս�(�H�l�o��(���3���:��p|�t8��h��G�����U������D֫�j2J�y�~�)���/���2�2 �'*�?��h]e�y�����h�C%
��&[�t#~j�#�(��ryj��K�*c$RU�5��`�	`��֊�ٓ��N��dD�90�f p#�p�6`�Yp�D�>V�A�ʡ�#JY�T)��ï��̩FK��{��W�;~ㆂN��4��¯��=�$���{QLn0��	s�vO��[a6@�3�C"w�<e3�2�����O�Eܭ,	F�y��󞱂M��8�f{�D�Q��i�5���,�vQ�P�d6(�QF�ؿ��.�0(G�0����1�F��~�x߽T����/
cy4�K�:2�]��,�CZr���0Π(�m�w[���'I��<&�*������~@.�9
P�-���`��-��[�?m_y\v���:����'����]�<�걶6�dt���O9{7k"2m`�Q����ه���KҶ>�K3����.E&�uY��:�˔��x� ?�Y�e[u�V�B�i69���}���g~�JDfYy�m}�~��~<����7���a� /��*Z38��0{�c����˜I��nj��u���|��Q�I���[���>�֣[�����v= xZ�nဖ�@�M��S�'Ex�-�w�?������f2|�0q	9��u�9�K���	.WnM_sz&�24*{k��7dݗ��+�#����|c0��Ne�Ch��|h��$V�x�w&���ش��%�r���R��S36�ߨ)�U���'��j�5�v)��.�J�줦�c�c�����x�|�ſ���A���	Σ�H��{:!�&~>]=�,H�����e,T�o�S�J`mc�YC�}d+����)�0'qA����M �����+f� ����{�k�>r�4�(�/�g��[���)c{����Ә^� �ɨC4��\�PEv���Վ�`�b�A�h�'��oS`�kp�%^��c
��+��g#�*)�PB#� )��.��"@q���~fh�:$@R�, ���'�6&��"e�O��Ų��ɛ��6���s�z3ԫ<�]jH�1l�0�K���*_�QDta���~m����dضl��@�x���T���Xh��h�.�:��	�.����(�� x�a*ΑKӕ�	�Ɛ ��cwB�9��e>^k����*4�m� ����ǐ{è"n-f�*Nm�Zh{K�*�W�#�5�����$zR!çF5�ou �S��4�Ex����)�Lu���#]opHfV���dN ���"v3�7����y�_��=��9�~J�9�n㇛�?�"�9u�2��^9IS�4I��Th���p���v�X���z�n�S���b~��i������9����d���+9�m�D�{>��@?���"p���-�9
�|˿dm��bȁ{��ЫKn�4���s�Xy ,��HEMS/���t�&a�B&�I+d�㬚���B�5�Z�;�t��]Jq��S��+����#rk�>��`���V��0��[\�ŅDU����]�.j��Iw��;��2�L�%Vi�qP+�����A.����s����}�I�ޥ�W��7B��e�z]w�"���R�Q��PJ��T0���F���f�?�4zgq��QjvQ�l���#��
���FP!�8�b�|���,�'��P�֕�*ױ��r⏩�s�י�!uI���ۓy�'k���%�;#�U
��!,Y��s1v��w6i65J��C�1s�B\ K�"��zّ���E�n�6Eg����h�4�,�2��>�ˣf����6&Y�W�e�RH���  <2zN��Ř��O.�RҕҪp�G�._�t4)s]1���1l�ジ�9�	��Sg�]�E8�wK��t�3@�:�?z�&Y#pn|kY�F�ܱ�_��队�;ݕ�B��џ����&^��[ޏn0����w�>��@���F};R�(�ƚ��SQ�2$͝��ӄˌ�6u$�����Wv ����.n
���%:�pҠ [��K���1W�XT�&H����]]y�|���eB�X��[g���ӔC�w���j�)؜��}�_��ޛb��������]�a�SB�<���'��Ҧ��8�;,�n��欿_6-���PL�|Ұ�~FW�(���G��}��͎�]�P�-�L~���8�0�i�.�B҉u���[�<��	�����Xh�qo��xl����u�RgE�W�I�_	���R���$]�?`�xh�$�Lq?3�?�Nl׷&^�z�xFz0
a�6���C�����qV6�"�h��rm���Н��ywE�V�P�w�+F�*�䜹�	�G{���۴��ײ��X~�~E&J�8�S�`�|1Zm�g
D��W�A�kCLk[�V�j��7��S��r��A�w�O�!Ɛ�کZ�v�Ή\�܂{���<���#FE:�3�q�/)��85�V*�a���->Bѹ9З25膆+cnY�t>�Nt77o�Y`��:}:�����Sg���]�����	$M)�/��8>�'H9`0��u�HMJ��\�J�&���nh�)*�y�� JL�N��C�E�sR��ש:�F��-g�}����Eƪ�gA��P�%� O�᢫Cڛ�y�0Z)P��\��y�zO%�q�/�q���?+*9k�l M����d7���+]4��`�)�f�Y�&���f�Zc�V�� U��І��	�G�m�wR�V��][���x�)�Z�Q�z{3N.-����K�.�Q{*�~�RA�hTX\�E�Q���h�/�̬ґ-��w�H���t�_���?l4o<~��x��T����R��-��@�'bE�OL>�bQ��9j $���>���'j��WNS���Տ�(,�dc��"I�JT�d	u�T�%�n�3~�i�rW<�Y$��R����C��ޏ�T�ɦ�-����_��.Q$��#dZcB;��]y�ū�S�����a�$A[�`�Z� 8]t�(��ޛ�ϔ��s�Jϥ'm�q�F�ƓG{ݍ�yy05%��!e�p��e��
�@ ��y��s�tt��$t�S��j��y�<1�3�I��y+*�-�)�e9������>��+�=� �ߍc��B�QxѨ3{/ʤ�b��P�/%k;���O-F�З}:�@iq��g��.�Y%�
�I;�X��m�&6mL>Z�1�ܭ�}����a��"o���f`n�;��>{����ɗ��SfC5�Htd�`�N�"U+5�H���[��u�m'&(��	uS��L�+P���[���0�[-�HV���Xhr|�@�6fk�����P�ާ������<?9�)�-���F�+ ��:�I��CߐX��Z��9��#�������#�Gp�p���[=�L�_��.ż�յ�k��!�����.��o�!$�F\i�:Y)?($稶��,��F��=o��i�Eo��k�D��lQ�ﶱ8A��4;�'Nw	���ǅ�?"����.
����Ͽ��A��M�C�#�13œz�������5�4%�d� n��/�o���#C���u
9�
�Qb��t�������Eo`�1���O��ԌJ�����!m���O�����5U�����>��c��ױ��u�g�.�[73v�V�,�~�ca�<�$L��Gښ�������� ��	�# M��� � 9�'a�2I�Ɂ);��ZZ�ԱX�.�:�E��7Th�<O]��>)��q�8��Ռ~�#-��_��c����3K�&�Z����iv		�����	ٓt��zɁ�9�#�}��J�>�&���� �?YF<�Hf��e���N���G`� %��0)v�O�%��]���,�����̔FD;��kCg�4�i)����ǘ��y:��н>q|�jϯ�P�K/=mY��U�_~:��E��d�*$G�C��,��+`><d�q����4�oVKBl;&���ۂ�5�����/$�ٔ�h�Q��;Fr�@5±4�~�P\�kwU�lY��5��\p{�ӻ@�L�P�ߐ����%����JC�W�8�޴��zS��y�"�g�Q�v��4��!��3C�ĵ,��L.H�d���T�y�����vy�U�$�$�J2�|���Wv9�?�f���(��dL�|�0���AV8����(�K�S�q��@�����3QU����pu��:C`��C�Rk7�� �4�����Yz���n��vu���Lnͪ�[���tY۶�7w 
~�66���Pǒ8�=M.�d�u�#��9���h�}�.� U�5��jQo�(j�]�r0�Q,�"���F�y컲j�����T6��,Z�������!���T[j4�c(3]�?�E���B��p�o鱵����m��Ly0%�tXTk��ȣ�e6�d��9e`�U��,�)z��x\�����rB��gC�>&*�����"��2oS,������ �����EG�����.�}�J��?r��\��(�]�^A��of9�q�[v)e���!��)�����*����w2	����)��\2�[�xR7���'ڶ�� ����I�P.˴�RR�I<5d�4�k�\�K�7��*jV�
=�bE/�{�XM����Yq=����Ԁ��9EQ��q�����P��Z��?�t���E(l8�C_����v��	�O�w�2I�j�ug:5%��w����T�*�yx6WK=�Ga�L��@�"u�.�^e�d�}�f�ǣ�9}+N�{a�#K��	6�8���vԲ945��`�[�cV����ӮS�(���(] �&�دҒ0>��j��G��^w�\΋WFٜ��Y�Xؖ*�;O����z�`L�krS�9�1Դ�\c?Ɉ� #	�}��C/Yg\�;�#)Wf�az���c%���⛏(����Ň@3����s@;���7Ph�?�Ɩ��Se�'?C{א1g�	70������(��1=��V�L�<��IP���;�>���aJ�|��.�J�T�ߛ^A�݉(tE#�I�ћY�/�a]�6l���{�Am��HL��'6���
�%��Ɋ�h,��޶����b��C�7�)� �	��q