XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x�
����ɲ��ˍ��Ǟ< �%CV�����iK��2�\�n=��˩�(��U���T�L kG5�R�ݙ��فf4��s��� ���Cyg�t{S���ӹo\������:�ՙ���`�m���}1�U�ߜ�LzQ��o�����Y?�-�.��A���(Y:����	��3��d�j.���-Ծ���c�b Yo	Z&xQ�6��.C�pG!pJ��W���Bn�aeՀAu7H4��^󻋞OY�baΡ#n{yQJV�$-����g�~TU�����p�^WV�霛�'�uV��K%f��FxL�so�۶n��nh�xv�G��}p��-:����@H���T)�n|�{��Kơ�U7>P(�;��q�r!KLÊ'Cv#����b��AF���8Aiը�����D8�LmU%2}��T޻�w�R�c����W�b;j
�.���[�����Kh�淲|�!�29mz�Lf	i�t]$� �'l�m��|�q�D�/����h/C��nӭ��	��-@��k����]�I��i����sIX7!�xD �ϚJ��"?�	YE(�� jv�����D�[�k��ne����W�CaѬ�Zsn~��;�m��h���ad%CB����4��e�Pȧ���&�Zj�n-DtQ�5`���HMh0�]<��q�y���Vi���C�b	����_�	;��ˆ��Q΂ �4��6a���[;zb����	%q�Qn���]W��8����%��V=�յ�>twSn�XlxVHYEB    38e2     fb0��ZN+ņ]�&{.u�Y�E�RK�[-��ԫ�m�C��H�L���Jթ�}�28y��\��XPڑh���p��	��m	�f;	�QSǨ��4��8�JÔ�LyrE�q�iΩ�x?4�4��w�nv�)f#ܱ�[�[Gy%'�'z����U`^�Li���3�3�INe[ң�&}Ȅ>H��y��;�	�o��y~G����om曹�
����j�� )�^"$T�MuL�wh�
�n�zh͕��dn�9$�H�kU�zF�=�D'E���@yqak���c��ȼ)�w��6~B�i68l�XQk+��':H��z3湥��7��l���b(q4�:�f�]7m>��4%����@yˀ� �Y�$*��,� �D�ӫqQk��҆EO�y0�/-��	�7���[�4 ��{�G�,�Lݷ��eߘ�x� �dK�/Egߩ���K����@��OD#���'q�Zua��� `�5��M"*�j3#�G�����h,b����C��*j~5�c��d�6��T�p�ZᏖu����:�~-�i�����B *��W�Xֈ��H�w���eO��6%p3���[��a=����g�F�:��vL?ʾ�!���@���#��Ν���`ٳ�/��y�Jv7g�	H�Zh��>3�>e�}��{�H��^�L^���D�j@/��5��Crʢ�R�V雄ŎT�s�a�zo�,��g��Zk�XOz<C�tD�h�l��p��)�54�C�)�%��\���ezREum���+���`�2�mn�Ϸ��6���s;B���1���2���:��T#��"Q3�N����U|@,�j���1��o1$��O�" ﱸF]��*6�m�f��1�vO��s��eO��G=���E/wcx��XB��Ko��-�Y�g�+�ps�6iA�ȷ�9�"B3zH�5%�\�t�'�G�P���Ć[́�J@ت|��u�X��>���mJ��"�n�G�na�;�a�:����������yc��1~r�2�٧v��L��O�����/�TG��S#'�|ģ`�i]�-�&o� ���2���Ԛ���+��_� �赜j��V��_�D���c<viL1�Dȅ�2z��`/w�E�j�cLޅ���^H��?�o~}JU�=�����k7ˆ�7C�Β���H	y���EE�s�{�����(��']�cm�Q��\I9>;�l�$w~!�/�4����s�h��q����CSs�B���SL�t�ޗ[�ӆ��߱���N2����I~���>�ڵ
KdؿTv��Q�,� ��.��<?}�ߋ�h+Q툏�BZ;�uR!�	Jc�5o��	��5)}2\�=�����"M���{M0�A�L�[�d�#�G��~�}�G*A�����:4Y^�Pe�p�Q���*{i�+�ʩZ��6�nZOڋޔGf�FS�����T��q�܀�"%��L������H#��D{N�L��p�0I
��#�v�u;��4j/B��Ő]F�6�#W�~��>�%߸ �� �b�%v֨�/L_�a���\��_�zS�'�3%�����V����К��"���T^mBB�T�j��S�F�ɐ��a��"�Ւ�LL[f-"�6a?&M�X�m)ܽ��-Ύ}���?��"AH�$�T4Έ����vߧU�D[��C�d����-N jɋ�o�-���|~ �"U"������1�̠��0�4�KJ������\��R�g�C'���>�t���A���C7�s+9\U���~�'���_����1,z1�_m�T���|�j!ո`�u���P���G���|A}�5��髃��Y�ʴJ�(@��V�ET͊�J.��1��Tcٱ!a�W��|L7��b�رkn<4�Q�$���n¸^�*�c,
�(*�g��~/�w�A�{��3p�
<����t�xcm��w�։�z\�K�X������W�s��ъ��Q�����Z%�X~%��<��H�DLf��6��t�oK���Uپ��_:nt��b~��N������>B0��D�i_7
���C�Tn�¾��Քc�ns��I.k٠e��~�g�����V�J��*0��=�zKw�&��QU��bE\IW���Gb#1+���\A5�9��u���'\�{(|�`+%��Q/%�{�\Z�J&m����/�&|e���Iͣ�!�Y�Zx�[d����>w�<��|� ���BL�:�b��}hf��B����lLϯ�#����ɈЅ�މ���{:>������1�=f��uE��b�z-�3���3.Ыg��G3��a>\�29��v7�gN�Xf��Rꬬ�ј&7�E������Y�s��]���Οݺ�ۏ�g�)�v�$�/��=b4ڄ�C����8G]��؂�&�"!S\��`����f�����Xr;���KB��7�v��x��oS���L����Z��F{E�i�X��Qa�)[��	F2���g�:��#]^�hG��G,�q,���S�`�0���$X��k]q���؇ `[���@+���E?:~A��1���#�p!���=@��jfYn���y�փ:��2=��!����Nj���Ѐ@}؃1x<F��߾ڜ�1i|�N�Ywm���ǀ0�~��>��h�s�l𰟛\�;���,���#�Qĩe6� 2�X'��pޠ�< ������[��`'(A"����Bc���|͊3����p0:�����&��(����w�y�i�3��s��+̷�u����� �n�r��%�#W�_/� �;����Qܝ���{1ɪ�c2���-Pyp//�� R�UB��7	ߵE�C}J��mh!���(^=�v��T�t��r>��IY���>ʷ�U��Ӯz���cp�	�����?H������0��ؒ�B���i2����SXK��4�25�u�d���l�����w/dc�4g���e�8�˛������KT�D��N�A��`&(p�wʢ���� y=C�������]j�@���B�!�Z�'d��f��a���ۚ�MI%��?�n��-gd��cP:��Й-`}�6�j:��{�a����j	���{�5��(aa�����*<�	6$��?���[e˧�������Q��tui��6�7��~s[�q�� 0����~TуK�r2��K����Ū��s�)��)�ĥ��l���l�p�o'9 L4p@WE�`>F�˻HS����b�2�L��p����q�9���q��|�簣����g�t�Cd� ���L�U��c��n��j���������[���1
��W�	��=� d���w��SӢ�FO���Ojln�f�|r��&q؉�q.Z��3��+/բ6�N���$��wK���F�W�A�`V#�d�}X��\!L�AJ�3ᝏ�;m ٪�&����ij�����.�
�RM b�I�-f�_���kN˰K p_UccIa�yf`bk�&�wAn���~] C9�����!4X��)����Ĉ�څ}ꐛE�_�{�Rƪ9�}9*��$�)�P����=�	����!E�o�I�	��m%<�5G�7�!�8�Ͱ�N�����h�f�� J!��Z�L���3��p�XKWF�@���G���7$�����E�`�Q��+�7P�m�\�F͂��|Ctc?I�����(�@������0���FH��#��.\˳-��ݵy
��N�u��eG,�s�Ǿ?^B�_@/._� ��s���w�b�QAaݘ9}r���<����l�5����K��'�  �?x������<?���ԁ�v����X����b�r�Ѯ�Zv,�1�`4�̲�,��G��p2�M�=6�/�������'����3�.��
����tva�