XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B=f�(OG�v��buc�>���-�?	�1���&��k�ǁ�wß%�D�������o\��>���I/8s��F���V���2��F�����x�/:����v�׺Tڭ��R0v3=�r�����87P�\�{��Kn��>q_6���0����@_�|e��N���ow��A�����{SNg�<��s�P�J�E����uש�LR
�y��"�.���w����+P@j7��r���C�7Ɠ%�R�g۸T�4�zC�l>-�ܓF�P���3����-z�tx:�i�n+Z>�;��ӑ^�ս��%��%؟�;���K��y�9>�W�o)�P4q�I �-�a?�N�eQ,��-!��T굸vC�eƻ�C�RA�]|�Z����g���q�2%M%���b�h�K���Ź�G�^�C��k�^�`���&~����|H�1l.�*3����#�S{��1A�]n��1�=���J@8�1��#O�im��O�H�V�U������z����v0��<�����o�~|���]�e�j\b�DRg!�c�%!n�2!-'�#��\���b�1r;�1ͣ7��kAjs��ɑ'w��&�\�BQ�ϐ�[��i@vH����XӋ�����0�S�Z��d�ɧ�}{	��K�7�J"��(x�ӄ�)ȋ�3��� QD���观�}$O��88C�5����ZښJ����ØYƊ3����-�&�� ���])����ݍ7;�n���*����@΍
��1��n��f��.XlxVHYEB    47d1     e90���9��bw	(tO��E�	�;~�5�_Z�sw�G��l~^�l��|4T�|A�v�HQU����M��N�ٟ��GKNp����=Z���p��nT��51�n3�Ɗ�R�6�F�Z��n��䶏�i���Ĕa�-S�1�bť���/ �]`���勖t�+vEE<~�{�P�&h�m�
��sx����t��\��p�>]o� ���l� L9�N��>�V�`�r��i�IR+Ee_�@J���l/V�9�_���et��벚*��'վcJX1?�(��8_,[R
}[i�:f��K�%\�%�7$e�tw�����ס�ϳt�0+�~��
��T��Yr�4*���3z�ⱶz�	�p͓L���@�2M	�+FQ��>F�g�A���8��ç��������wPJ�/���v8��4԰+�Y�� �(\���z�?�K��$ e��:^\��<O|��b|�a��r#��u[�q�u�^���rXx�ݸ�:�� [�K�`�O�,7�T�%Y��sJ�(�(&�+Ej��#��X��������ȯ?���:�S�͊)}���ܝ�c_�&d��f!,V_2"�h]�E�rD������yԙ�K�Ct��A��B�?���$��yV�y��%�ĿWX�s2�����#ٱ����z^~���c����m�>֠k�������%���\f>0�A\�"Q�M�fֲ	}p�"�)k�l�!�'�'�#t��U��ctg�C�������|�S�ѯ� H��h2V��Y��.�9ZqK�:-Hq�������l�~/P_���G�3Ή�ȫ��Im���9�ւ* $�\  h���V��������:��~��1g���4�֖P�d�'(���6�����5��2��ڹ[MY���7ǚXR$��^}u�\�v���+Q��ʹ����kUx)q�j�"��Ȝ�t��Xś�x��U��*���Z���2�ȎV�ړ&s�<�]�}�|R�z���;�$��쨻�EĀ�_�Ii�(� 
�n`�H����i��X624R�-ߐ��e��4�!IQ3����K�L�px�V��Qj���R�!I�yu<R`Ӕ�?��ٕ9eh�� ]tX��2��� Nh�C�s��8�=�9��������Z_ͦ�P���r)xc��������Zj��ʒk���T=0�|���C�Q}M�3�w(H����Fu��o]����WشT��KD�(���X��{���uhѳ������kp��&�M��7t��yV�T)dN�M���.���Ih[f�1{Q���b���������� 9(�=t�xb��=a��7���e���0v�OZSj�t��<��~�Y����bnչ���Je�[�9,�d7]����4L}+�s,�gW�i��b��KvR��c���d�,MI$�� ��Y�&T��M�'���J�A�&0ԭ����JV�n��)Ue���i:�6+Q�H�j��c���׷�F��	���2��n?%�,>XsK,qne�=G:���բ z8q���*#Tz������(���igaA"YT����K�� ���+���7���F�6}��-��\b��[ Ж��%y�܅�"&�c�o��dW�&.4�fWׇ��z4����p�4D�p���8<�Q�Q���r+����	�ef�a+W�d"�_�U͉E j�s�3�Bu�egZ𻑽���%�]�op��uʨc}C� �AJbE+]���3�χO>��]�%vT��7�J�X7
�W���M(y�T�8�me�{�鉭Z���v�P��x���ٻ'Io�W^ǯ�]�P�G|��]'��b��~7�n������m?[�h@��{��K��m����A�����f�i��7_��lZ{��.��O7)�no@����\l u"ܱ���S��T"�Vb)����x���E�T#E@��W��?y{�m�V�J��R�N0:�Lģa����(�d�R6 {n��w������N�E�f���������gTWj�`�أ���T׷�BЉyݭ-�	����LV�����)��:��i:��,�2tA����iG#G%D�f��M���ʻb�a�@�eu4a��me]��>������Gu�'K�A�:o�'m�i;���XE�o#�+��Y�Dm9�'9��s��`�'�&'p��z�X�Ћn���F����d`I�泽��tI�4#�h������$WF5M,A��3���ݳRRi�F��J��O�d�����M�����.~��܋^�q@���ܷt�gW�S8���Ӫ@	(Ũ.7c*��R���D�0�+W��5��%���|v㛖��[m����YB ��?D�b�*d�1h`�t?f��vݹ�e�� ك
��R�Ɂ����HG����I���d��_�:;�j;+�.�sP0�[�p����nƀI)K��!�a�]< �3u�[�8Ӳu�#��o�$Z��3��|���+�R��W P�H�ZNaD�ep���~�b���hH!�R���*1���bȚ��G�$��yV�C������߅0�l��b:�ko�I%�$�=�G�������8k!#���xf���5�� 1gvv'��§�b.�D��;�d�*��ym����˜c3���a%
��=+eX���ց���u$�]O~'�`�˪��n�:h��w^�!qҍ��t���d�$�8*�cn�	�~�J*�z�S�8w��:�;��c
�A5/8����l8\��Y� ����璮�D+�[s-u	��5�G�S�,Q|��v
��������6��a(u��;��$:�b�6���L:it���J~�*Z��J:F�����r���hHo��ԭ�_>�e�RE<�=��������nվ��y��UMr�!I�&�7R`��?T�Y�h!�,$��N�Dze�������*D#+-�4}h/�z ��)-������E*k�}1�s4T���D��,#uuu�K�#�A�2��*��ﻨ�_3Hv�@Ӥ�1�=�?���0���Np��\'+�߱슂��%_�j��Ճ,�j��H������ |k��L�T�A�s�<_>o{��c���@}6�_�2B���?N��L��� pJ�4�1��
�����s�v3���B�~��n���������᪰�a������N1�Ti�]��e�!5.}���aO�*H,H���w����iT���M���R}B��ٖ?�Yht�w�����;.Xp����Og�@o����*���B�Ƽ��0�A�����IDE ��@7jk�SO����[h!�Z����|�s�A��(Je�Zn���&�9@�&��R @@�I4�&H��r/���:������᡽;���#�ڜ��0�&�2�l���ګE0�/��)� K�(�_-���,M^�uFmhn� ����	��e��0gm^NCޫW�o'>$�?��N�E�ό���U�Wv{�g��o2}�/�Ь�,u�W��y�"($0'����by��#�k�[f�9; ��8|e�Q�fL
~����Ա�����~"�4��s��/�}��M ��-��y��kv��Y�k�(�us,��#�.���ږ8�V�ZL�o��sTbҬ-������A�'�KeR����̤���|��o�ح���;�