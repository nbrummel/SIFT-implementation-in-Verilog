XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������;zY�z�gj�8m���OP�Z���H9�a/���#�F��9���E`�<��#���^�F���[���]�����A�X��b�`�1����Gn��	��]/@�އlT`�k�;���}�x�$�w0X��tP�&8~U���#&��ʸ2�M��b��=*��m�T_
��Y����M?�i.�&2�/F�'$�׬��^Z�%ZU~��r��@�ES��x=��ҙ^}Ѥ]�a���\E&���[Pi�(
��J1ɟ8{�v �u~>c�=	|��|��t���s�Wu��Z���g��s�ϢN_~�'�$:E�RU���k��b�z�/ǁ�80�>���$kK��j��dq0����݋���
$ۜq)y����0&�mbu�Z�:~���<P'x���Ҟ��y����8<遁 Gi ��y�0<v�����E`����RX}у̳$J��%�s���XJ&��s���2�\��fA7����*P<G�2<���(�54�JԲ��CLax�R��2c�49��/~��º��IVfmD4��&f���2+���l��x�/��D��)���2���l�)5�He!�Pg�
d��ڞ +�Ax'um8�\KLNS�=iq!�Р#�K:��j钘X^B̅7��|��A�K�x�$O@Hċ��Oo�f���$f�V:s4���s�>U��:Xх@��yՍ�[҄�K9�Pf3�����O������R<���
Sw�[o���1�XlxVHYEB    fa00    2240���%�z��t��Nǯ��'�������G��(kQ���M �n&'��M(��=|������N��P�	�=�K����ԛ�ٖd:w/'��愀�蜆�@�A�uv��M�[�i��z_��w��B�jZ)��'��)��4!e2���j��}m����Zг ��7��'
H��B�-_x�[4� ��K}=vF+v��	�"�\x���ŀqz[\-z�d�|�J�P�̸���1L��:[�"��2Y��X�[L�����jG`6��[ՠkY��`����`��G
������f��5.hb�+
1��(��h����m| z��ȱ0�A��x���ѵGH�}ϸ��V�;P(xƸ8
���&*�bc`��x�&h��m>�kl�N�j5����vFiH�A�I��o&���wd������p#�RԾ�X&�L������])��`�Bq֔��U���v�.�-7"IY�*D�4*`� [��h��@�c"�-���0�rM�F�����U��W:.R���fb��V��ƻq�F�C�+L�K��H�+5&�"GԾw̌u�z���_L�W��<զ[�r=�z,�X���)��'�n�XU�/3���`���xb�l�4����dW	r��LTС;�~�z�"9��*���2��@�k�H�$�|��M?�;ػ.��I��2 ��`���9��Ր�XO�;��&R[z��ˇ�3ta����<�WwS���
!�V������n�=�ck���gh��f���+�	J@jG�U
d Z8(ϻ�;U�[K�Տ|dN9G���RUv-M~�0�'
����n�8����y,�@�$I�:�-�}8&�����|�W��za ��Z�2���c3���5��^�ɂ*��z���e��;y=�Ƌ�<318CIEMc����ھ�E<`&r��*��YB��f#����(��njެ=�e ��iCY�D��kJ��V�midg�ad<D��i�
#%�p�Z��!G�X~%�:���a��b���O��P7{���Ջw1��H�"��H��۩(2�>@��ZT�&�������Y�$��A0���ycq5�|����o
Z��@۹4��z�MƷ��r�� �p���&�S�~���+��p@���ރ�I_�����"���&�dE�'^v�i�r�g�M���[B��q��&�5�t[)0pR�2|87��1�QI����SN��@9��R���	�1���1b�$R�����^�)L����܏:���,�+ł\	��"C�kH���_��p|^�K�������'h˼���)
ijqp��_�8)�65��7��?��T��#�z]&t���� ��vZ����L.��8k������*7d��=�B�
V�
K�	�+�a���w�ݗ��*����abxn�CΆ�P��£\�	n����J9g��v��7�%p3���5��f��B��J��~a�����d5��<x�k/�y� K\��c����s�7�N[��P�Z�+��_���<�ϰ�*��v}/u���!���]jP���P(�U�/*� +G��sA�}W[�]"ߐG��^�q@<���`�Ĝ�:�/�tL��C�������
$#��zZ+���a?�鰡p܌$P/��z�o8#��B���~���] 2�nq��IDf�c���q�2� /��+2AIjN�����1�N�P���0A�z4j��33\�$���X&�����¹�������nb�~�d58(�%�,l�^��h��*�P�nB	���ͽѶ_5n� D����O�$'1�G"���WW}��Z�]�4ӻB6��^�-�փn)��a���eϏw��-��O+}v���]\"ԟ4�*����<"��#�'�Al�$B�E����@�EfPT�H���S潐�n���|b�!{�����f:�.a)$�`o�����VCl"܋��XL�P���� ���������i&�T�|�'0<�ɦm���&�l]?�89r٤i�re0^pT'�׭}舒	�5�o� �3N��=���G9f<�ѓ�6A���Qd��?�ME�	������Y���g]L�'q��/��t��-%<�cBm[�n��_��;�,v�M<�r�������H�$��e7���B6���,�W�m�K4Ss�M?	�__��-����^�'�3(<p��� ����/�XM��O��"��ɋ��k���J`l�/h��p�[��}A&�ضj��2������+-V
TrD_��?�C��<�;!`3�X�v�O���mI��%\y}
l*�R2�[3f`K<;B�`�� +����N� 	ʍ=�-�ޤ� �& ����&��;��o��,�݅��vǍ�� [r��oҰ,�{����WW�&u�$��K��6%׳�� 	�B%�@,ʛ�;%�h��#�q�\9N��X [���DPw��23��K-aV
��j$p<�x���<�y��l��zH'v�����ހf���6���_`��a�J����E���F7�KD��F)������}GZ��{�����20�toa)%YX�5�Fn�qhfM�V�\l5-s_n���_�F?BG��q�\N�Z�(+f{	K�ӷZF�8K��7��o�\c��M���|��i�z�ԵA��M��&+^>��	/P�Ju��ct��7ՈK'7Nz��t����2#hi,����6�vIF:�וE����K�o@?�}�VN�Z[��5BZ�R7�A����C@���!oW����Ma���Ϻ��wCvO*�B�1%���k��ѝ�����c��4+]~q����{0[��Q�'& hĝ�ȸOq:Q���"��oU�5si�g�0r���Y2zV�Xs�rR[���:���,5�_S�4ղ� ;V�����(�����\�w�~�-(��_4��TS�yx|���]���f�G�Ԡ,�7����L�����wQ���ʻ���4���U��3u+E|�s_M��i�-Б/��{4�J� ����븬B|h�!��[8��Għ���b�����9����Ύ;�{Un�*��W����Ӆ�פ�k	u&�t�����L]�/D�����w�Q5�e���ü ���Q�� 0jnH���5U���=��ˊ��{O����Ά4���Չ�'�Q��ۃ�������5��׌|��)��&�,����嚶9�0���,�V����Cٲ��V��MR�Y�֪o��/��\F�6�ڎ|��l�4���ӄ����$��]�����aZ�����6��֩��;�ig?��ftml�Õ�FM�+\A2^gh��}=��p��7�qr�ޤ�	5
(�֔JGy" �݀��j�{X+V���'�O�V��i+Rc�˭E&V��R#8�k����]�q�a�]w;G%b�({uʪ��x����8F�_.p,� ۡ�x����)�~�B�P���4w4��7��m�@0i׆HE�!l���l?��$��E���Ԇc�2�鏢"E���jי{�VFՁC�2��5��CخўY�mUl50�nړ�W)�Tl����W��P�F=3hj˗mq�~�~�h��b�Z�&� ����μ�؛�=��.�0VB�~_ ��Kֿ�89UeL��p�-�xy{�ui0@�� ��VZ{��J��S�b	�txD����~V?�$c̶NXt�`�1�~ VL��6��^��x����i�����w%� 4�v�xF��
a{��^���ma�wER�2<M��V�|��Y�汶.����TL>��[�g����72h��>��s�-¼]��ת(˩I�����=�}��^�TH�/z�3�2���)˦Do����lX�φ�9IT���0׽M%�ՊA��x�7�K��;�Ld�Q,�[ZʸxGa�<���y����B��%yM��i
�pbAޞ�յ��]�������EZmQ�J Plq���ǆ��z����c�[R���mIv~o�H��iagT+H�;������H2L�w��Ʌ�=��W����t�3�{*��c�k�a�.��^��ˤ�`��˟��?A��+AZ'`�-��;����D����I��`T�r@��SF�t��{;̜�*_p��TG��S,Q5g�U�>0"����ܰQ�-��+�� ���bx���LȲ=H�V&��S��3˯DN�%���.��rN��'�AMF���=�5�Y�ϼ]��/�K�z���D0��'�2C~>����Zsu#v�]n�u�ޛ|�t}�/�Yړr(���a��6-1����c;�$"I>���D1����u�����*�q��_!�Q	��Y�U6���P�d��C1����O��'>�Uu�l���aRA'��7�q4��pe]kQ�N):�����2B��dL������j}���a{ܢ�j���k��:ȋ�_��	;�w�Su{���{S^�p�<������IL���N��*��ͫ��e�;8-?
�H����%�ȇ�֔�^��.r�0�f�����bk���I��U�+Rl�36�`Rx��e�N:��/��|�����":q*ՄΒ��W��v��봹�0?�@�,�3M�Ө�K����zIR��kq����A�+2fWX_Ɉ&~�kz��CČT��\E$c�F��yż��FJC_�I��#����E|����+�3�Rmh�k�ۉ� K�(����ʾ��]IX?��\�dzZw.j��:pPpB1ؘ��s��yLr�4Ӄ���ns:�o�3�*W�9df�����$D+�+B�������悎�K�/R�IB��#&�)u����@�Y,����S���-�a۫���O
�P�l��) kc� �BѨG�/jV����m��1(��L'�_�*�C�"MV���ThO'��@ QHMuI��zjxx������5wA#�;���Ƣ�	D��qhA1�/ӎ ��x����sĆ���v���U���,��������Y$�W�lgwe祼�>݉��.h��"�L� ��@9Wg�J7��4��V҃,e�����Z>k���$��.\�Ŵ��w쀛���e�AKD��"	�-c*Oǃ�Gz=�\¨z����9����pA�4�������,?o�H{ZbB���#_p���g�N��<����0���1��
sXc��u�i%&�>����䎯�e�&�����߄�S��W«�����4'�_yI��E��!�[���hU&Un���J.�4ԕ��lp?�r�ʭ�,�Y.��E�Qŷ:�,|@S��E@BF>�6����I��(���H��@ƛa[͙���웗��Y Կ�e�YC�*(��#���d֚�K' �j| W�I��i��;?���
x�l��M���%����/I,��+N(k?@�)��Z��蚰��I����[�vWpQ���7����u��
a�,3?o)��ͺeŹn�:��C�(��Q��@ۖc}%���$�fю�~	%�H�����1u���H9@�G��M��<�x2ѬxI��]d�p�m#77���(��������]j���_x�� �6P҃;"��ħ[-�����E��.?I/��I;,E0�X�v�f�̜¹��
�l "��v���h�Kh����!�6E]r$m����pb.��z�9��5o\�ov�*5G:�;I�8���h�-�̮�t �:�@�d�w@���C_`1⹀"l-���M���'Ğw��22�\���ƨ�B�஍ �N5͘\��]�;76�6����L����a����e�8��d[7�*�U�K��3h�a伡@�d�m}I4c%�
`SuS�Ư'����rفѨQ�� ���*O��Q�L�"���t'�+�/�W Ab�JA�<���ű�:�d�,���Fz'4򦢚�q���伟��#�ג���.{���� 򽅚y2Ϣ�#���q�>J��$sbAG F\��pBr�4\2��z�[<��k�:�����B<(Hy�lN���P	M��B+RIfO$��_��4O����M�u�y
3m.S2n�<�,�.��ls�6����|���\PD&�:�<�j� ����[��,��N3����N�+%C��fG�2x�c���.�@8V���ǧ�<LYc�&��*|l�;�sB�F�BDas����]��0cb�7���f�w���`6_�b~:ci*oѮ��%n�O�JU���@?ma(3,�n>1�hv��o�+�wL����g�����y��Ӌ<��Jl���w%��J��t��2���5D��G�׃V���px|��"/�9��VMD���r�4�c{�N+�kO�O�O�4�,�iQ�4d*�!'���@��2����ht+�D! ���=��(c�w����#��ЫKt�F��\��Y|6&c���1̾�]L-�S�蛩�ch��a��6(�m�pݢ�F��Łc=�W����v������}�����`�4�\�"-O0�6~�p(�z�m��A�����a�����W���V_R��M��8p[,-Y8��9hM2	�q�nƶ*z�_��B�#��ؤ�Y0���i��t��;�:*'���H_nV*��<��$� �ĝ������^�J5jg=�I��M�xpظg؆�{)<N�`M�6�������E��<:��Tzl\&P7��q_��*���Z��
G�?VFD���{�׾|�r��!H�
 ]��o� �қ�{��	«��vk�`��F$)<W�����H�LD���NM�&��r�����3�|���>��'�Kf1�Z
U٢�N�9���'�܉�<�R�Mmt�AJ��ҷ$9���<͔x:�9]�il�����UU�	;�7&)8b�C(h�%�qgcT3k@�� �B���VE���i���t���P�Y�(߯fJe�2��bM:h�X���ϝ	>��R���i�V\*Z��U��g|����m��p�l�h/9L����W��w�J��|��7y�<BS�M��2Scl�Z� C�i��,�n>��aDK��a��ؤ�f�h��s����֧{>�M$�h�EC^#�t��QQx=x��x�  �����b����--َ"���7`T�`�>C8��2�T�'WTG�#!�mAJ"ŏ����A�%?��n��LD��S�b���F��Z絩b#�vLE�D4e(A�i��S����_��v.X�\lbZ�s�.7y݁w�[���6W����y���5n�\J����~ik���Q@��GQ�W�^c�
}<����+R#�@�+���+�:`J�N��-�g��/�$�R>�p��G�d�G%����,3
#��o_J��E}G�93�V����ʂ���%@ra$�u>����=s7E�C����}�Qr��>lѢq�m`��i#����L�m`��J���6���[�oT�n:5��#vF6��P.����Xr7s�3�5�~Mg�4�pTr�R��!��HF�f�Z���0���������
����UM=HJmQ�2_�mse:1ѕ�%U	p�~�/�Xot��n�6*�O�HdVq��5����->�j��u�'�4�`����b�~���}��0����)k6:�1ɝo2�;ep��x
e�W�$đb�3n�{P�ܹ�`����_0��)d��N:Y��G���i^@>F���yr�p���h�jb����M�F�ƭ���h;a��Q$��-��s�JЕ���|�:e'�=�!A6�%`5�l��@���B�||
af+NSi��`���8�I�@Ȕ��!,�������1�D�x�9�pƇ{�t9�?��l8�t`�C}�toY,�x�N�����H�O�s�/�O���3A��$��0b/�2Q���.+������"�YH$F)~q~V��l)��5O[E��#;tЀ�;����E|�˄<���7FC���K��N�����ո�3g��B�2q�/=7Gj�QJ	��J:1�:�VL�*�@���BY50e�
 #��ăF��rvc"`evx�}a���f x��	���>T���؎S�x��߿�f,�h���Ei7T���FV��<����Cvĕ�Ԉ�D�p�����+S��̴���s��e�6�����E]��&�a[k������-����$^�{���K#3�����!���X�X���'F��Jb
+�`!�;[B5) �!�>3T��L"��r)%�E�	�hm#?[ȇP�u�Z'"`1x;�x4ٯ�2N��u��L��ڰ����y� �"�|�z ��$ ��ɽ��e$,�ՏrȘ�#+�X&�_f��$�+P��3$���~b ���7gſ�υf�B�M�,�96.�,�����w��B���+��G��M@�^��L����VcR�U_Y���׋���j;�\rk�1u���vF!�ɫ�՚i}ZlQjY�dI�����i�� �˓w�����$m��Cj�~W��@��8�A�5er_��X�_i+"�]K4J�E+v\�x���<M��¾h��n�s����nŊ?Z��;fj��_T�v�+����g���[d����b<?`�=��c��!��"�5����$i' =�A��:��3��T�x4�15�6���j&g�O���L�^̯��~�|���.r�J�}��|B)�� ���L��H���K�W�7�)FR�XlxVHYEB    6682     5d0�ς%$'�[~s���"�~�^����f�"~m+���sD1@�G0>������f)���s������O�6�Rfy�[�P��6V�����x�Jx��EI�n���ٜ*�\`�̋��"i��B�Ny<��#��FA�Rɇkͫ�Y���is���F`��or	I�*`m����G��Z2�7�.g(@YR�� '��*;X>���`����N�f��":N��5邍�LL�o�K� �#m��V&�R�~�!]��wwʗ���rs������-E]i^�j�ɹ�t�G���R\)�(_���r�*x=�h"�]�i[;H���y�&Z���k�c(0IY���aNIﰕ`�P�r��?YR�U�o���(�GJ:O����U��]���6$c�6�R�''���������b��:�aY�4��Ӓ��Q��9�vq�w�:�E{�~O�Oh]"���j>�c�3|�C�I5������˙�f�@��ȩ�$�^��@��7#?��^�0���Up0}?��=h�zȄs����}Y�B���(�<u�h)���q��k�<G7��D2���{�na�h��/}��d�qaݤ��b���m�џvM��	�A~�^y����갏�����W=9��K� �g�H
_��5�w�y�41u��5uaE<�	�a5&$��0.�%{��@_phޣ���R�U���Kl8㒉����ݘ
�f,�)�3���_6-u�շ.]�*�h��
iUO����_P�A/Ҁ1���μ�4�OӱH;�@�;�i�Ҕ�  ��o�I-�odCC}��B�����	�~L�Ue_<6G��z#��#i,[���O$��.c�㬡wj����\�Y�w���0��L�K���S�:9����������6K���ƺ�ܘ�t
A	Eu�����\QZ���-�[N��Y�R(T�~w}DD�[��0�{�����S��Ѿ� �o2<���~�Je&�ius��u���YP����D�;���R�І�!�2�G�9���z�<1�=de�vЁ@�9���L<Si�iy��SP��xZc�4�����9y5��dZ���׋.��i ��!�@���L�j�H�!�ى*����T�2I;��_Wk���<ǵbǵ��@g��/�=��2�	�쪭B��Px�rK7�������/vח�y��2��?����F��H�K�qr�,�p7�#�<���s�����R?ț�%��~*�a�rzbIS��)�w��9��2���2;�Pr%���5��Vݤ�b6���xGy�C`�CK��rE�U�����/�)��l�V����g��[���E�#��%P��\=CT����z���W����g���!i94_�s�+O6�A�������f��;�O��E�X�1�����#Ŕ�°����.��"���9�r�zx���/ �7�Կك�%;��L)x,x�by`�+��P|׳�}��