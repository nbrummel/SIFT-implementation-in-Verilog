XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����D[^ot<J�fk��))>v���+��_��:���%L&C��mm3�����V����_d2�L�=�փ�$a^[����@ؓ;����7��n -������S�D�[��{���(<��3y�f�Q a�9&��Ǣk�H:a�CH����E��G�y c5���V��])�aC�fn�-�ܜ������.@9L@덽�Q��j�-� j'�-ń;��	s_0���Qq2D���ڱD`�_ޣ!��,z0����;\&uo(0�b�[HE�]%PBY�y��n�0\+�*���|R� ѿ!�3�)��������;��=/�_*#�����q�T�W;cz�gO9�H���2po���G�$/#�����[d��'�%u��D��T�O'�w�;F �s(��^{u �MXv}�`����bS�/�TХ��V��0���F�&b�\�Z(:��=B��,�=b��:v�Gس�����Z�.����+"�l6��d_�{����M�W��d@б!Z�<\�����H��|E)5�.�;cX��_�ߌE���>�7=�@-]��Ѐ�p&�0��u4igg?D���(rL=��� y���N���p��q�*���YU"�f���3��nĬ<K��'х�E�kv\eW���É/���e�c�����~���8�k�wy�'6/���Bt�y�ȼA?�w?''�:]�G=���͞���g�R�{�{/�+����ԇ3d7 �?��mԳę�B�K�iN��x]w[�/XlxVHYEB    32e2     b70�۹����"A�^Ҳ
A(Cup�����^����y��Deϐ.�~��>l���4�x��[uɶ���W��2}�} [$�o��ef�&k(� ZA ���l}��]�M��,/(!�a;W=����4M��}'�qp��k��0����,�����鯛]7�WD��Rq�z#��ꙻ�wM�pvF[ ҝ��u�\�j<�/N�9�/ژ��z�Q�b>i��:B���_��E"�,�{��Ώj�d�4���E�؊��6!�|��1\\o`�A���z�ߩhx�H�(�^/R�ak��:s�@2�mn�nv8��4{W0���6�J-CǇ���m���_͍�r*��!v�hb�N�G�3���� �u�c-$_��������:n�u�(�q�1�Kv�g.R�MǓ8'P�r2bԈL�����hy���=��"-R�������0zL'2��������bZM,����:��I�'^�x�7�)��KO�zt 'sk�1:�|D�9\��ێՐ�2��@��a�K(:��I�� �=V6;(�f��I���(N���e8�r^)���X+6�}71��V��R��MK Ӡ��M��l��$�uNs�VV�*�ءaS�9�y;��\y�7&@g3=ܾ�0��kC�U�R��ݵ/�"S�/���z�z9Ϫa�	���૎��?\�g��C���8��C���ԦS�˔巣�e4%�H�����JI�* X���T�?wX���Oʂ������TY��"#�&E9�u�b�$/g!�.�vI�@�-'FܨE�/]�1̛��F� �{�\Y� uM��0	�t]��$ذ/7�!'��w{HcbgO����eO�J7�H�����sʶ�K���E��-��NR��eY��V�
���\�o�,N�+�5bR�"�+���>�Mn�o��(P��[�+oƷ�-��.sō �K����93[�	�5������/���&G�cҍ�[�AGA�5$���Ғ��Ÿ�4����mm���S4ҕ�`XL��P�h�f�e"	���>�l�1#_3;����[���va��p#����ͻ��S����V��QxJ������`F\]!�T��$=�F�����*^� ��\<���+�jD�jXE��Q1�p����[�CB;�Y쵙�pS�t[ol�rL7$Ci{�nWɮ��Zk��{�-,��I��*dS곩)�)}���	�t(���s{?��$��h� U0pqW�%�M��������w��xj<��W@�$��IuC�_M���CX�5{�=z��q;�\uY���=?�����x���#����PC��*`t�}�.{���о��1W�c��My��P��=�j��P���}����~ӊ��HR�G��bQr���]RN��2&x3������:����|�Fi���Ѿ!�͚Tȑ�4v����z��E<�W~�?�C��6�����䰽0�m��Pr��s�e�����?}� �Τl0�.	��G����;�/,;���MG�HLҨٰ4�}���>�J���꙲7��n@ꔪno�r-XgS9w@Y�u6��0�s�nE��u��:�|�"2��8��[�Ȧ�t��*����S�Ij
δ�2����OsT�S�!��sz�͑���D�Wz
\<����f�B�z��`0Θ�M�nO	!���P"X�SJD����H���O��U�Wg���x�ЕT����ϲ%���64𿍴NJ�Za�y��q� ߈����>�y蕂#R2P��%�	�Ԙ�a�P^&
{����,�k)�\or��������f���C
��"�T���Ǚ��M%̉h} ��L�s��F�f ;�7��w[����p����ߕ��ݒW�/2�C��G+V�Z��sY�,c���~ذϩO����l����xfٶ ���_���=�� ��a�32,\?���L3RV��C@95ؕJ��uW�/���kB�r{���Rq�����
���Kʒ�C��3�V�ү�j9��B׭;ܞw셸�'�B ���Y|�H�be�"�5?2KجZ�NC�QG�7��>��aA���zS�m�	�)`~�sā���*Og�dt?E:jw�eo�^��ԵZ��G�7:kK?�͍҃v�B�cv83�=�lZ��#E�T�	�2\�갪�,�@�B"~�Xy	 ��
��7V{f�+XH]��4&T�Ə�h˶�j\��{=?$Ec�����^�rӆf�6���+�^�����+��Ru�ʚ9j�B)���-:��|��0J��;��ꢕ��s�U� #��[��U�ʣN1��-��,�$�8��^��R�JŇ��d[������7�c�;���hԎ�l��2J0� �# �֥���D��������w2�Կ��c��.����S͐�����	(B��}	l�!1ՔEe���0�����O������۾K������p��el�Z#wah�HO�t�@�"Q����2�q��ޗJ2��FZ�ԍ�R�2���j(GA=C"Y�%����&q~��= ����Y��|���4e��?����t^��M%�ʕ����B1�� P3��a*�Y.�����c�Qf�^�N3���iH��/��N�$*����iXt�X��c �0}P�+S�*V�~r�k����(�.~�S�OeM�ɤ܃���� �"4��Qݓ������	�ph��$���̥����f�D��4�Y�"/�]Ȼ�ϗW�XF� ��40����P��i?L���5�p ���KV�!�J�wI��!���u�/yrE�8�I]���
Hs�%k. ���>�����J��X�ސ�pj-@�[5*��A,·_y����������n�JHN�Äy�!�X����d�x"��Lx