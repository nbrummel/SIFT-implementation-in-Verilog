XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ot�&ݓz:q6��ݗDDС¦�D�{�J�D�%�X�8���Ck�d"�"��)�t�VԼ߻S�q�9:G�ue��
��ʄ�0�_��L:$��y��MP�R�� ş�Ĥ�F�ե� �+X\ђ��G�
^��-ŷ	<�g�ه����J�P�8kQ$]Y��y��.F��D�~���d��"����O�sGg��^�;�b�z�ft���o��=���R��B\��FfQ�¡x~���<^!��[��,e���#����j�/����a��������7Y��_�t�� �{6׵��v�3c���	�/�0�
��d��Ɏc'��9�K��gN1f��K�dܣlY�VR(zÌ~�<���*�R4�2��~8��NZ��E�d��z��艀�k�q���-]os<V����_�PL'aqL/��c �
c��Q���2k���xY���%i�@���{� ��!CEjiԍ_���W�\��N�r*��a�c��,����'3�3$8���q|�Ǭ4Tj����oe��)�͙G�r�<�4Z 1�\h��=-롮J�Ĥ���;lL��[v�&ɫ��4R�,�
o���]6�׹����G�K+}ô�L�n�k)?�`�5�0��rr������$��Fk��j�	�|����n���ś���ݹT�Kss�����m��"P�riY 1f�\<u`����p�R��X��-$A�������5�~-�k�-ȡ9����U!���&���C�F���jI`��F^�%���%�4ZKXlxVHYEB    1c45     9505e!:��=+ݕV���a�%��)a4��Wm[bD����m=���LcQ���"k�{�K:�ܼ`���h�#[�^�8&�8`/��Y�J����f ou={ �?�MFOXŏ���Bފ�
�`#����#�3r�
n��___O_�*����o���N\�Aw�+��󫝃�R��?d�ٜ�f�}}�M���aqaQ��Y�%A~l�
�5���W�V����i�5�P����[�����\�sh�fԀ9��)/W�!�R�2,��)P�ґ8�L�;{��0�G��k�w
�2�0�&)��i��灻�Z��eU�\`�_�4W������Q�����7w��4y�C�9�&u$9�h��/��1D����d6z���(m�*�K�'�n��#���cu_�k�*���8��ٿ��ob���0���8,�"p?�.J=J3Ȱ����%6-!"��Q��fH�kU5�t1�N�ײo�A�%Y��k���㔮�����+� G�&�W��6{�T��ZO��D���qJ���ZY�ӹ��{�t�ڲ�C�5�id�O�9�sS�F�6}4�֏>�J��YFlKgW��F�@�n� �����l���ի���4�`��C�߂ѿvJ;���0m�����������$ΘS�\
Z���tz�6��\|[���յ��y]��"ֶ�a3�F�����k0�``uVq�H({�#�����}���,$�ZB�p��{y���]O�\6׌c�H}��L8~ǶnlGʷ���v�-��AWo;��{w�8=	x��iBJ�f�K� �x������W��G�vv��P�\�~�m���,�$�~�����t4+������X�:{r|�a��im6=�Jp���n�P'����Hᒿx�}BEx��NU�F��y5}�E�Ö��)�ojҡ-QA*�J�j��a�왹���[j��\0��S�S��`�3�����v�`�R�7�nGcp�[�AB�̟��9�o���0F7b�)�s@b�:ش�M���G��}��)�>=~&���/��K���/X����-�rg�. V��d~22Nq<F�̚��l�9��}5��a�����{�`�HW��b�s��k�8�v��5Ne���*�\�a����~���0�!�c�C��H��IN&/��h���ug�D����i[���d6dt�bh��L;���#�[J�1:�H��벃ʯH}�m|�8��@A/}��-^�s��2 �w�:]*���,��t��I�z�1�D��U��VzI��Q�95��[h3�'!�L!�(��DDL�.c+�����#�>�9�Ѵ�7A����zТw�~|����헡qtLV����4r��B�~)�"Ok�����̅R���QTB�}�}E�����)_h�1jp1��cߺ��B
h�}�C�p�엊���Bg� 2���%�Y�����q̺0��I�R.��}��Ye)����5L�7T���g���ߺ����F�F� 4[����۴'��$�'����^׊��Ĭ����]��j����b:��ꈏ̥�%�K!�0�ny�E�g�ȽqT��#�#����(����>�Z�(�Z��]x�wQ�h�ws���	[�	T�����hwcR#�,����N����G�uF�4?�&@�����?�3b"��S�c��,>;�S���v@n�&��$U_1 9�{7Æ��l��!���%a��^{k���Q�������������k�7;����/��kx��kf=�X2��_�&����S���hL� zWR���J����!Ӧ�l�
��FW��_T�꛻ơ3�?�ͦ�%�w`�T��O-��� �l�;�_�+�j7�7�Q������YIׁ�e�H�ܽ���$���j��fvl\򴓘��ϴ��U֥��S��Z�t@��,���^��}�&�`O��X�}n�U8&��7�u~}O�0?��w�ێZm`Y]|���7@�����$��^�E�{�	�뤏��z�s1��N^���Q'*�:�!B�9oN�&3h�K����� ��d��S@�*��y^�7쿩����p�gl�	q]�Ƅ($6-�G��t�	6����W;"$t�֐6�s����b���g��&[�u��b�@#4��@�ǰ�TV�G{�ieR����ǲ ���y�(��.���H}�u!f%�:!�����h��e����vB]X#����Jnӥ?ٔ! �pU�U��uC�`.5>��HL��o���-,.9xn��qT_ ۼ@��a��Z�^s ��:O���K�� X�\��/��] ��o������ݏ�w9Rd��S��03Q*svp6۳+�Ǖ$���kx�