XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���e�e͆�sT��$�~�]o�+|D����m �Ƕ�l�(���hyKVm���%$ �N���/���ڙ�~r��n�E�/]\i ���~{��k���c�J���}����s�B�2�5['=E/�5��m��=5����%l���i&5�4<��ɞ�׹~�uD��֥�7�<JX^z���XVP�<)s�/%7~�l2�4�c޷_r��0�=�o�a>�\���w��\���.�yVz�4k@�[@?	��$�ǟ�8�����F�e���[�x�33�m�Z�!�p{�3��rժ8�G9��/���i��%oj��9�On8R��aU�xT{��_���^x'Be�"�o��j�ܑwx����d/�2�k'ݻX��lrΒL������ܑE�	)�Ja��TR�p�.�^�%W*��iY+�ʪ)�BnOl�?3�6�����zt�Rb�f\���K��X�C��]�Q�(b��؎����d�m;ah�n�#���Yz�`W���ڵ�6�T�9&#�K	 � _%�\�(nx�ᚓs��9��U��F�uL(�| &7�;�Y�b�X��w�%�h��^��ݹq[��}���p&������ԾX~��h-PA;��xlZ����g�Nt
�Pb�iFƵ�pҿ�>2`��Ʀc���*��`��hhԆJI=m�8v^QC��A�3;et���N~ufqk�la���hO�QY5A��Ɖy�2��EU�����tx��P��֊|�q�;�\uo�`�Y�"Ro@)�XlxVHYEB    67d5    1150�4�y�c���Q4^(�S�8�������f&�1�}��Xf�5&^�3(�0��v�+�d����[7����ڴ�G��}%�?<?���D������.5�ἦ#�f1��lQ���lْ�%�^LiB����)'����B����/Ns�YPߥ� x�*���u�$f��Ha��O�
I����'W�DC���+�8��8��KM��Nv�_�����eP�!O�bNd��X�c�ǫg\�W��	_xc��12��]��yo�Z�dW��h�C%ֲ,��I�T[�F�����+�c�^� A�L���|L��+@����tv?6��� ��_�<�u�_�K��ȿ	Ӕ�,:T 2"]7�jb��FDs�w��wDG
%��� X�Q�Q�@
��b�Z��`������3Y��]��r�lktd��LP�ǅ���Ϸ�a
2unbA;Z�2jj��g��7���P�H7�84Wۺ|����$���SL5ՎQn���t?h�5��vnD���3|�01�=�H]�蚀���L��X~a���^�5�xֶ��l@�;f��؆�Oa���@��=m�v�-�.�*>�k�QN*/5:M��KQg�Ҝ�S����5
g0ߦ��ZWd ���p�̐O;�{6~�V�n?���N��2�����h�"�2E��h�a9K<��������{��w,'�}��I�=���7ϋ`]���e=H�٥���pR�S�Q���z���
~L�k��'߷��4�5�8��5TPs(���X}��,�B�mS�+7��k0T!^ϑ)��mS�ߚ��1�_��f;Z��+��a�
��h�����g���]TXAp)�=��	���t��C�� �{5I;�:F��Ib��<��~,�����ҴTr��wb�2!xD��FL� �mj�|�!y.Q*�l�c�4S4��|/5/;Փ��g÷��w�|��^&�Z5�}C��7�a��{x�+��i�7�,ފ�i�L�2��3<�2��t��يB���_j�-���B���f4�UEK��\&�pE\��ܵ�Ń(���_�3�'�j&�t�]�YE�
ш��)�.��kt�sn_~g�_��'�����]��� ���Blb��W��f�((lD�k0�ʷ>��Ci���^88����7{iˏ	�Gs�~j�Уo�%J�*�o�L�x����F��5���,� u��]v435�a�݈|yϢ���ϊ�n�������-�~����ǐ`2l!��fA���sl7��P'W���^�ڈ��E[���ڋ�)���]�"�+�����Ff�M�� '8B�=��z���|2��J�N�1�}GA�t.�v��n@3�Hx�F9��*�����ɔP�=ܮ =h��k��0������AF�� 7����kU�@�;#X��?nIv��+�~�.Z�����5A#Y���ňơ�3|�W{yuw�� ���Y�ڣ?��\���8� �-�M�g�}#p��K�)6\opc�jǉ����=~��q��<}צ#'�ĝI�e�d���r�Y��h�l��_|M���:8r �2��,eBX�V�
$��Z6�A�BF�tG/h�Z}�#_<�"كgh��)�VF�91���vz����)㯭�=�� �����nuH��/M�JK��2�n�?�7D�\uE�ߺ�H�u�.*�zO�$���&�,���2����κwt�]J&��C�y�ʂa7���(Zғ�GFՖ��ʌ��� �_R���ǻ3�TQ���-�;��qdf[l��C-Dɋ�cJ��W�]��~
�@���;T�}�����{�����s�OH��E�OL�Ǜ28�/xa�������5m}S�wV��O"�ק^uB�7ǽ�D1k..���s�f�$���gzV�����wMt��W� �z�6��I7"|��v�WE�>OQx���LۍӔ�})����q�́4�A�G�ѽ J;R0�U�S���u�mrQ��WHM�tx��h1�#I�k�=#����g� ��ɷ�|(��ø�0�^Ze_�o���[ˍÃ��h���	�#S�G���mC��e��Ŧ$ "}!�`HV<� �^M���]q"R���fQc��&׀���/�?��-۬�Ϋ��[����H-���S��눭�];0��]l�"!֚�Ar�MtJ�jQ���H�0�q�1����7���J��D� @9j�(A{n5�$�JAH&R|v��v�3�K,;\L6A�j� ���%�C�G�������Š���k��\�7�1��CvI[��xu�A2��r�}���:��=�Rٙ�t7
����Tp�8��^Y��4	x��\�]�Q �<��ԩ(����� �/WԷ�V��������h`��%R��Ou�:'y��Kі���:���Q:J�o:��9����p�~n��������p����a�U��X�����㖲Z��|1�,3�:�~{3. T�bX�Lװu��`[̖)^!2����[]G�H
I"��!���`;����N��M��U�d��Q��]�����9�ܤ�(��_�DE����gͧF뜝���ye��Q�U�[,U��x!4�L4������M�"=���^<�|��;���0СS���N��.!'������šh����!�A��hs����+���<�YT���b��R������6��HB���R�v����z:G�*�dǱ��sE����S�	�r�x]\��l��ʖ��2\�J3�v�x����v�;�U��Q��a"��"�z�z3��N@l��g��Q�J�12�,��l̚��S�f�����$�m�⹐�Z%Ōw�����Y�D0���c��,G�O�؉o0���o��Ɉ
���n�"�-��`�Xy��2�U�3��P&�vE݀<���5��evV{2����aY4ʇ�]�F���џ@ �(���6Q��fl	s���1)e�o6�����]��y�/Ů���V�"1e�?��t�ԍr���b!{Z7��P��b�WҾ3Vj@P�#�dbs�y��e��ri�'4w�u���C�R�ڕHǥ�q�ݩ]�S�S��Ku�(��6�Z�i9X�ˤ������O�:���w����K�Ky[U�t�L9�w����R4��?2y��R2��o�&�E߅�@��<o�g}��os�A�V�t �gp��{�t��h)��Kl��r��\/�}��)I��"�v�4K��nxENIܯ~mq�7���SVE-p#`Һ�"�"��[&@�o��3?M&ItD���̓LذL`��et�R�b�%"�����a5�\���[�r"����������<�'V6SJ錼5�w?.Q��5�zdac8�'߶�+Jǧ�j����)��S��O�W:0C����au���?{�㰶W���XY��͢�;q��t�L�8e���Z��B\�*���G#��4��n��7��V��K�c�H$�|96�XK�=�R4���#�-E��(��0��K6��*��z�<����v���K�t���-�GS3
9�[]k�y��zbj��'�HT��~�δ��_�BthV����Drba@e�s��{B�3)ڴ��<��_hc7��✦��|ŖՐ>S�A�y��T�ܢsc�b����4����JO)os(��P�	���4EQ@��a������"Z�=���l�j�Q��2�π].{Z�2��S�3���l5n�eC��~�
8<�����^�������.�4Lg�#��1�.���� �ZP�X��
<W��i�4����j@ �nT���aw=zx��?,ڌ�7r��E�AJ����*t%ޢ�����0���<HOD�g�� x���.���+o�:��{k��y��wu��"��!�Cj"�a6ϑ�P�z�Yb2��"�$�E���X��8��\е���(�d���`�=X!���yJק����w�\5n��_�&阖�뜉r��L]����|@��<݅�>꒪���{^&��q��p&�\"���{�7�kD=&Áq=~�98�s;(����d���?�F'�����U��w���ߋ��8�?�_�ߠ?�>��'t��� ��[M�gQ�vc��f@/�1��C�Gj�0d/^����+��G ��li���������p��%T(�����_j� ,���M�ެo�
2��S �kXy�.=�۵�:�G������Q�@R��]^;Jdߧ:���u��P������?6P���>rˣ����fcZ�o���:9w=4C��T���Sظ������Ѯvu!�O��JY��v�:J|4�Ǯ���W>0B��!	�wɯ�$���3�5h-U4a�����