XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H#4�������l�gp,��%C/�'�5��V�+f6���Y'����|�K�%�.`�س������Xf�O�!��d<`��U|���/�jXh����k�ל�ʕΨ��N���Õ?�A���yT6�]+4��I����lf�p稆N�����p�b�W~WJ��FDr	4ӣ�R�f�{#�� ���>�!�ZB0�����R-V���$�d#���#Qy���F������W�ke��yܑ�(����ތ����[�J���J����Jj��6H�%C01!%��a*��z�j�R| �E�� �/ޛ/U�M�<�ٮ=y��Hr�e�%��|;�>S�Y��k3S�R��/�q�T��qi�D�>�����w�ǖ��TP7+ԉ��Ωo���l�6����NC7.ةHi`iA�~.�i_{\����)�b�O-�+q�Ѽдꂬr4�$^W6&�5���R�s0�+�Ge�5��n�&JU���G��TF��4X�z����&j`h`����3J���5��1�P����Č>�y/�C�xNF� ��1m X��9���j�/��k����a����Û�����P��SJt��ч\�}�	� ��֔�LQ/�i��3�[����`�l*"��>k���	�`9�w��#�ٕ9�=h���7j�Q#�s޹��%~!�&A"�cS�Mģ��ql��Q��\�
-� �	�ը/MVܒ�ٸ�8�4'�ؠ��ss6���R���B��Ξ�J9���`XlxVHYEB    2f9f     c60������م�b�~d�ɫr�@�4�8�hz�����C37�c43�|���y�>o��{��d-��$U��B2��ƭ�It�r!D���zx%�Yǃ�ْE�����u� ?	qHf���>�z1����V�I���Vf���[��S����l�7J� 4�J?$	~�ɑİC8��5��M���t���U�&��ȳe5�߄P���+�Ii�ʶE���mA~�҃3tۺk�Ó�wo�,�����)���v�uK��=�!�l	Ӛ�����3��^Ur��*KV�Y�i�pÉW�%��(9���E���U���]�I�\3����Ŗ�&2g���}� �.��i�W�mX���ZH	�e�	�:	u_���Щ���,Z���u�"�\�X[���۷Z�I:)c,CbBZ�ʲ=�[�[,�ׂ�"�����iKc�wkd�J�/�*�i�A�T%���k�ke�ݶM�y�f�aa˲f��
�Ճ��h3Y]��v�WI޸J�� )����
�R}��Ǧ=p�����:��XE�{�Y�#�z�������%舛̟�=@�_t�J|�q~/ܛ.n�΃}+ى��r��^��2��B�\k�moh�H��	e�h�b�#F�ߗ~����'[�;��)�٥���`�����U�Sc��S�
F�T�u���Ǹ�`tp���u���w��޻-(�w�^��ȗ3-��b�l��\�i'����,�ۀV�����w(��C��}#3w�D��������1�������j��U�ۃ�6���g�?3gѮ-a��[
Q^����z��g��Nak�M���fyOL��X?����x�c�0�{�����o�h��H��L1�E0o =�ZxYh�d�}&l�)���\h����[A�m@���2�+Q5
O�N�CJ5GH��;bS��g���,��:-W#;�%}+�4ob,����"WI)����,�?�/������,�u�dr�L'Gj#	b]N7�����:ɜ�/ǁ$r_b�Nv
5
���$�ho������r>��@n	�x�Nv�0���{-��on-�i��h�&�G4�����"�� ��;�2�#֗HTT聀��j����f������0h�����5b�*�"9e˄c�v#�\�X].E�}%f�'����	`kțH����I8GݵU_"�s�������D��������D�z�#��h�a�=F�r��Q�Ò�7���#��G�:��>OJ����)��?dH�����cR��WW�)�ӑ��	�����y�� ���U��P.�V�������4�8����>�<ܹS.����g�%��2gm�"Hԍ��g<)��EQʮ�~�,�/d���)f�����q����ȯ��vP�I�E�M���O�y���Y��T_=1���@N`D�k1
�ݤ�g(?�8"wԩ_)'�:oK��I���0+O07N\�3�@�`
�(��J�L��9���5͟��2��& ��С&��yz�
�����]�f�lq��%��U�<k�q��P�����M5����8�1h4��e�mvQ_k%�R������0��D~>F�$�*U��f�}��9%�ƙ�&	��K��bZ�K�+��=#7�k����� (U;���|R�i7 ��P���B0%B�_?��G��π���e�W¸��������dM�x[
_�Q����f�wQ��غ���bR�l؆\����%�me�;�د�Β��ڑ�σAJ��3(�W%�s�>I�U=D0Dׄ�d/c�t��B�5Tƣ�g�C~@o�ķ5W3��Z�P-c�F���V���09M2���2첉ݡؾ��ӕqm
zC�"�puz�>��}A.�SN���h�t���i7�Y��ϧ�G�&���!i�qp������v��F���R)�Z5����
����i� �=�7��8�b/��boz�3$a�%Sls���0�� 	n	fF��U�������(Xßz�k����A��]�<��{&��㕬�G1�N3��H�l��-�����8�B�F8���G�~�o0M��J�KX����w��z�Nm�HQ�0KN�+�3�d�1����B�t`�ĝ�#e	��O^Z	�������U�
=�qt�g�f\]L�y�Ҟ�DQ��O�Bz�@�{E{
aܭM��Iv�O���]����!����ۧ���?�����b��3D�G00Y/����VctFǊ�2VWM׊V������ �s�:tpAw��r{����V�4���."f����S��G����"�Zi/����Up	�>Y�����4�7��Ǒ�v������e�'1ft�2^�~�d�d��`J�C�|�À�N,�2f��G�7�0�4��QOvp�9l�{��2�	�jC9��	���;�]n�n#z36��p��@���?�rTV�$t<���,B3-�@�*V���D���H~TW1G�	��J�7�gC��K7'@�k����]
���Zq%��G��g9���@��~�ꢳ!XoEZ���3v��]����v�L��c�0��z�˛%�2O�-sNKz�~��s���i0|	Rz9�� �fH�<����^|�|�._V^1�����3�8l*ePqεi����d�Г���).ځ�c�b�^Ֆ�r4,Y�aɚ�<n���U1�_�k�lO�p~�aq�B7S�<�Z S����o:@�k_�My���k :4l*�G���m=�"���O���5_��3����޸m�"��07�����l3Tt����� 9����/`�Ұ���6a���j::�y���>dp���j�q�ǺF��x9��#d�/eKv�����D��ܬ�C��RUr��б��I4�3�oմ����!@q���3�Ҍ�[����}�z"ʖ*�� ��^�4[�<`u@闰Lx���Z������p���Zıg{P}����㩼��iD^�j�`�D5�}_w��A��i��.A�(�ϗ�=H\��҅����5L�+�.H
9�3����7&�{�߰;%n*-{}=����c��ǅ�Wr�e4�	��zl�V9�F�*��R�e}�������O����J9�Kv�(�]�6Ŧ��˙����+���