XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����M�
����b��A�ܾ�yS��8�J�]��Z�(Q?re����T���b4��]ʦ�K�<nd�E��i���LL� ?�0!]L���6<ܻ5�OZA����L�1ߛ����En�������>������S?��ʲ�I,�Yn�床��s�H�����_�j8��t�F��k�I=����$�9�(�0��Ŵ������!��X���3�#G1���w1��X��mMr,����Ԑ��LH��Qih��A��u�?���������<�OBٟ���J����h.hG�L\��SmV8���1�*�g�QGO��-:�]�zM�ʋ�^Tc����΃�����l�A��`hwA�����̱��8J'��#�P�xy^IO���<��w>}�SSo tUiV�5��&�R^�o��(��t�"����q �Dd� ��j�lV��Lp�Bh�K� �ܚ�c!��[Ng�Z&�����&"*�z�y�LPN�������0�����ʹOu w�����&nyh�g����:T��@#��J���EQLo�Ά�몮�gjZ�QL��>X�TT����H�C��m�)��y�%��@HQ�AEH�|~f�������>�#C� /��O,*�kܝ��8��O�QF9)=�9]���xc�a�Y�o� p��V"�� W���P|��!sG�=�ިUQ}\P�n}�%̩E ��^Y��i�v�35��B��D47du(\��M�	���n���z~�ޮ��l�,�*��-Q�XlxVHYEB    9732    14d0]��S�<M{�	��0���O2M�!y곃�u��k��ȎuLD�1��3��p$��[$er<3Z65|�/�ٻ|3h[GS������*��{5��`d<bu�0Ĥu��9�olkq
��w�����?d"D�Cޓ���� 7J����[i?s8�E)o
��@�G�ň�o��Dd�[_�T�h�
�`�|k&�j�n[��q�]�:U�cr�?I�4��%N;�Ż��Lo2�-�ҟ�B۝C'����YW:�[��[��x�KY��M��4|]�.HH
�н�N <�f�#��ږ��@���לd�M��o+ސ�i\ad187F��Kn ���o,kn�����_"�3�9��Xh9Zʚ)o�B�\�$�ć�s]�4�&b���Nv����TI�Y�b65�M�n���)fR[N�9���Z$�|�:+�g�I6�Fb��h
O��#�!��:Ӝ��hzC�"��~LKx6���V�Od2n+�T#R�!@��N�3���m��2�/�F�r/�$0�h�Φ�
n4k:��Pa�z�Pmx`aєe�ԃ(3
X�V�@n�jV��<�2��y͎'O�HtjϞ�7(�'��X���R��IY��̔lЅ�S����q�A��՛���������	�N_AV��"���&f'�)Ʌ5�09�E�Aե�ݔ�"'�w|+�^]�-�20�z�@�B|BsՌQbEgڌڿR%�V�����J1�PA�4U�-Z@��x����3%G ��ߨt��.���K���<k*�Nkou�f��1�ү1�q���w��\�r|�=�'O�eAu�mx_cX��疿��]�
�cZ&?hS�.��1��7��{\K�B/k�����e>1 od�rv�(^[���l��N���G���2�:�Z�\n�owl������H�VT��&�ᚁ�"��Óu$w"X7 ,}!�"@�W��a��t<�J���9��O;����y0�ַI�C=G�X�C�l��!����3�������R��Ҵ%ni՞�j|3�X~�
Œ�=R0�����~�A2�<�X����:Ϙ��?�a��`�{Z�Y��}!5h��E5I;e���s9���&��t�{�ږh�QYy��L��Љ��_R��UW~��l���0v|X��#���@��/y�&��UK�H�:=d�D@0v�O���:ʑ���Fs��+��ɡ����ι�b����'���j ����r����	�]JP�-A9�A�^U/�"āy��=9ҷ�(�x���>�$�l%�u>j�<�:��-l$�m����oQ��7�Kuwzd�C��f�&���k��b.�%{yg��V�U��ݐj��4������b���Z��Z��*�b�|�-V����Cp5|���o��]FJ��ǻ�V�GT�u7=�l�MY�в>�v��s�����n_�I��ɹ���E��;�Ȱ�q��oa?���ct�g��lo�������6'xIʊn��Z�5�n`���x+p��V
{�`��5�fyd�pQ���P�'Z	�vru��OaV-2bֱ�F�zx^x%�lzv�zw�/�|�H(��ֲ6��iq��c�6��� ?}tlj�/X��]&C���qDG+��Z��г� \e����� !��������{ �W`��N_�H�!�)�R��sF�ו�7{3!U4aY[���!
g�eH��[}N�j�;��>g���[���h�SZA�"3���р���ֹ�r|Q�
(�Jt�w,PNI+��z�*�0<j��L$2$��V�ӧ伛�u�6������{{�9y����D�fշ�f���Uu��]XK���Q�
�GYIj �E�&��������m��w@�=�y{��4]����t,MK�]��2��3>b
g��n�Ŷ��,.��G�9/��C2����O���:���;H<j����d�����D��Չ�V���g����6���)'U��#5�/���}X��3��k�@ �@�?��|��o0/���Y
�R�����|F����ƍ'�ĵ,��Ix��Pe�\��ZA6��Tl�4�Gx*��hԦ�0r,۹ֵZΧ�w�s�M���r	�4���߂��Me'�
�T15�\�ٓ,e</g
�|N�-��3����2�(�]����hI&�*�����a��j�CH
�R�W���d\6�e�w�����K�I�)�|�O����G�����"�$l�d��dWT v�*vY<|�r���}eVQЎ�s����W��H얁VF��H<b�;K,���xu�����$I60����3t Ђd0
o�`���H�AF`F�y�h�1�R{i�8Vr���t��QLP)���vZ�^{��r�7�0�߰��L�o�{ �2"Yz�VH>��ğJ�D���+�f (�V��8�i���,�J��xnw������/��S�ny*C�җ��cLr���+y�	�$#�6Yn8�0]�-<͘%���M`H*m*d�^��\$��!�����[n�:� �r����[��L�U�΅m�m%�8�	ނ�biy*΅�`t.�{e>V�<���@<��8;3!h|�ݮ8�{�X�@�M�O�k��Ԥ;}T<����,��9�n��� �n����c��-1�A*V���0u�]uu����|�p�*�H,Ez��.�7���b t��<�.�/&���O��9���]D�8����p�]Rl4��w/|���G��5��v���OA5�3��h�c�l\��>qx4	�Hc�d�:�	�u"Y;K����cŘZت���MP�S�E��f�s�t4hW��5Hx�w�p�h����.:���S$*���TX��xo���s�G?�ih�šp�Ν�-�ŕtʜ���mc�괍�u/r�j	o}C]홙B=��d��m!�,f����e���px^����Z�˱fm\�fM��^�7C㈬v��?�kɣ�3T'�0��Y��9v���5oD΄��C��ͼ9��dxy`",0��;!ͷ7�����F��KJ�n���FQ"���QGcF����e��� ��a?߃��m�K�O�,����ϥ��*�`����dc�]	ҲV��/(���;s�'�z�*�%L�����ۣ�F�F.����
��T��;~�oeR��-Pm)O�5�B�t��Yg�=83w��V�7��f��mj����m�K��UU ��"Sl:p��Шm�s��<���y8<�A�8E�bƿ�[ng���3���>���L��Đ�a�U�s���7�������,�E��eL%���/Ͻ/=S��:�[��T�;=�?�t���h^��v*�5�Q�e����hˡ8̽����]�M�9Cv�wo�k1"�\4:��s�~��z�H�EX���<0�9px���m�T��W�s_ޠ�-�DP�����Es��Ģ�}�_�:7^n��T�@W+!��%����������h)X�+��횟wik�RŸ;����?9F�������X!�.�I��y����i�_�3�����P�c%�TǨ_&�S��~tX�/C�vN��}��1�'ʗ[�!5��Lx<{V�+;��xN����zW}���/�Q$�x�F�hu)�<�>��ߛ��% �(˓�,u:Sm��6�N\H�僼�SR�Q���#�
�Rqkq ���{A�[m�� . *��%%���2E��t��K��?�#��\{�d#6�c������"ϑy�o��={|8�,���YH� r	%�N�V�o�JV4y�!el���gg�bJ�t�n����J��кw�r�����Z����X�WK��o>{�b�9TY�[S�N����'?�J��eAO�K����/%��)�k%D��a|S:��ۡ���*�T9�R�����5��;L�-��4�!B�j��%=Z�'F����x>%��`8�\��l�PPƄ���y�}"�nI��k	���ٖK��j��{�9����k�mGFW_�m��
z�<������� X�\	@Y�J�%�������{��dp�!��CW���ϲI�bC�z8̋=_��XNa�u������"��(�>;..&^��Ui�������qZ���ƕ�˞��|��z�����Z��CO���h�\*T	n�$�ZoGw�\i=�����}���%:��&g�>�U�OdUi�t����=0<�-��3=�u"��#�"2�c��]�92鐌:��=���oق����܇�� k��]����Du����������0��g�n�m�/�����?��s��H���]d[�&A���9V�]��#��6R9����#�e��J�sk2�b�NE��^(�w5c_�<�fGc�?d�eS�ʯA�C3�A�+5����CFb����G�e���W��_.k��hx�?;�������������;Һ�V��x���|!���<�?P�ɟ��y$F����U6����q_�C`u�ö�Hc�
���!�?`Ȗ��j)���6��r=����s�?�����|Z��Nf�y1���uH����e�������d�g��w͑�#����-?=�?\Q����+ւ�����A�f=g��ʦͬbs��(f�:���i��w9k�&j�}�<��Ό,S�r�m�h|�?��4&�Y�f�|��L��e>��ѷ��.��2_��nn�ƶW�`�Хd{t� L.&m��������~XV�#(��/|OpҖ]��d���S�Bآ��fiVyψF�9�Y��<����[CVѪ��}��� Kb�U��Y�K�9��!�.񷺽�N����o]H��\P��4K��4ӽ�hn_������` ��E\d�@@��RK/���e�"@���N�Ȝ>�������>�#���~��=�2�r�6�G	���U��ԍ-$��ydL3�]���5�UJ�؍]��Ug�( {��?W�$�����E��Ź�����,g��GED�:�.�_(�6wꟸ,$�cg`�	��~*��_�,ȨS1���`�\<͓�7/�6�Ӯ������Y<�XE#w�DX<��H崗g�,)�5��/1\�I7���W�o"�=�R�Tob�p0��_%W��ݞpF��f��XZ���g�t�gL���y�ډ�3����3�n+vx���i�G�Z�8SR�DcZ�6�`��wx�nd��뜀�</�c��N�c���Ơ#1C�HW�1�"���Z�ym	��z�fΦ�̶��a�§�XP�'3J�+�{y(GMm
�6W���]�/�oh�%�J�`�ˢI���݆ɢ�#