XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���>SR2+FZ�Ό�O����*7�D��p�Tf�V��������H��عo&o�F��N�Í����Q���ظ#jWU��G��Ύ*�@����tt(?ټ�x0m��������ь�PbM]4���[��*��Y���<iI�q���6�m=13�����I�Z�^xT�˘���Ĩy�&MKR�7�E�po2r+G� �`]��p�#~ |"	*�[^4�=,!J�.�'tM���K�V�>a�3f�W�@kSa:��ҵ�7ݩ<����#UV�<�?�F��5�Ly�MB������ܡx�M�~	#
�t(C�ꖋ�au��6�����u�m�c�Lo�'D��qآث$Tם�HyxM��I�Ӭu'����6�:tJ��Wە��2�@Е�_!�Ȍ
y۔�	z��"�A;ri�3�!�n	C���^��5BZ$`�oxF��%�Պ"_�r�~Z�m��ʉ��٣ݫ��:z�s��g��5���3h�o$tֱ=�Z�@�S	����ǿr?�{q��iޏ��5��3%3>2�\�h/x� j'�`zvݮ�7����Z�jpW� M�E���> ��	��<E0��7��t�-�Ի�;o���_�M��Gɏ�����jeju�%�(,-�0D5aOP��>��ؼ:Y�;k�·^��֨��$�/�9/�p�8��Os�h�L>5�����C9�+ZNŋ��#�W���x�26e˹�VMr�f�����x�7&�@Bl�z׮�"�*XlxVHYEB    130e     7a01�ۖ~r���y�wl�A����k�v��Q�c\�a_���q���Ĭ5����`��$;/,��ypṧK�їi�J#_~�!hdG7YmuEŘ�$�8q��N�Ru���ʋ����!��p�^G���m�^bV6e�2#��� �?�#@�Q_33&����>�[L���Ҟ��tt)�)��Q/��6�@r����m���&�/���Uԃ���$�vV��i��-(2qq��P�}0��Ұ|ࠇ7U��Ҍ2+��Gj��yXZXѴ4�y}�ß	�_�TX�����%I8'���� Z������ݦB������9�2�,��;#�L�Y�H+d}�e��O����K����FR���٤�5r��@^A�Ϗ���_����)J�:�yrL����\���]e�|��`����(��'Ԝc�Yw�4{��3��!@~0�w;��h�j�f��nY_>0as�k�|Z�]n'J��G�~��o�?�����w�8�ecKM�*���k>,~L��b����Ќ������z*)Nik���G�eYu?|���v��$��9]�W]N{LU�+�{M�or9a���	j�=>,0�P��c�"e�Y[ �<��W{�cJs�,�j��o��D�4\05�o���bXx��l6�e,tb�
%�4��������
뗣����Yϩ\��NBK��z�iM?F��X��k��.��u�dԙ֜�zy��(%����J{�ڱ�k��L$%TO�����P�IoQ�?��b+�/���V�NX�.|]���Y�$.�-G'7�Bp0�H`\-2u��XWP޿�N$^Č�y��@�nێ�9��Qr�r��[�`�w���_������7i^o���U|��{��'�ùɈs���ɁK�^�N�����l�{V7�~+@d�8�w�gs����|�]����B$����TV��w~��q�`#�]�J�[�&����q^>�e0ϝ���=��U�b1<�uǣ��S=��� �`z��i���u%\a���E4*��|��Xd �:-�I���6�B��Ǜ�B�r!��D)Ϲ��{.���1�]ԎJz(�)'��-S�`�_$��=�u{��{�>5p��S���~ݧ͆�4��΀̖��gų�>�������"�ż3̆R�C�B��	b�9�pZ����������5#?�h��Y8 ,�t�D�ޏnz̈́�}n8�\��F��gs���������kC�)"�ǒe�V2���^�(�G�v(\iSYay9F5�`��nE�䆎����P�����w�|�!�T��f>��7S���ܓ?�Y��H^��R��g�!�7�	��G�]��=Ӟ��������
#�'k#O�2��a:�����W���Z��i;�V�����D,��bL�̤M�7T��d+��QjI���<�Ǫ��_!��e{�y���$�A���՝K���eO���������)C|m1��-SC����Y��<��K�}X���ۮ��w~NM�_/Q��U�'SpQ��d)X�px�P�O�1t�-"�})�K��R�p�W��~�������k�bz�n��e�vl7f3+^�S��6��ln~<���+9���i{��<lÌ�w�F���,w b�P�.T�+qD�^!Pd��r�؈��B�΃B��|*k�I�͏l� �� n��jx�ݧet$
���5��h��M5����\���>�`�B��F7���t��a "U�IEY6-|���E.�q3J��B���l����i|l�֣���P{��p����&���ۊ��z��d8��L ���h%y��������׶ �!���e����ϼ�1vr_Pfw�l0��H8[��rIg"�~��c��by����p�A�q����UD-:�