XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���1�i��ez��hT��ңD����{$�L2�\7[���L��r��mtf�{��^)ģ��������M%H��w*m��B��`p�E<Kɩ�EM�Y�\@~�t܄�ܕ���4V:��5�m=��G�HΓ�8<����5�g�^���"a�\��|&B�>�A�q��!�y�ujJ*��0�*��ǈ�v�P�Ȧ1��i7�W|�!�M�6��hnV{��S9�J�F_��8@1�u��ߨ�e!��wx��0F�
лWa�w��5�Z��'��H���4"o��û�ϙ�T��PXѿ��)&+=A�����+�.�az٧�Ki��e�<�ç��-J	Lo{���[߭��	�/3K�t�'��� ���X�J���_p�T��X�m���J1��Z���c�=/��'K���G�4�Tfqh�[����k���ٯp�ß���h�)�Ә]*�G�AT�
��m
��y�����t���ݡgU��d��NA�\���a�.4Mf��rBϽo��8��������v624��J�j�۷�N�y�BN�d��Ue�ꐪ�����n��U��`��܀4�S�[���hZ�A�^HIqB
������pĭ�,\+o^�Ȭ*��0z�'I� ���Y%�8�|����*�Ya��\�-���#�=ZN�a��5�o�ل||�bF����|Đ7�EfI±�L�'F��U?��ۖ�ް7JXǪ�<X��T����W(��TGU����TS���Bf��̷���{t���oO}XlxVHYEB    8e9e    1d40��|��I�U�~��ްz5�SL`�m|3��Zz��c;�E��xR��p�=�7����^�"�s��D����=4s�Q��L{�� ��(
;�z�e�$�>�����?;NGOB�|T��Sqޞɰ�� �M�|Z�-�C�|�-�Q8�4b�I�9	H;gI\�(�i�����S^����9�g�p�e����v��ף��H�.Ѳ��㰛P����7�Z��ZRƖ(�f]�XJFk}z`r�n�Y�=���Ss0�*�[���^A��V�F=�A��FBDC��j�I��W�?V�M��N�d��x���u��4ع�E��p�
������o�r�{��f�:.�V�7�62&Ί�4����d��p���^F�, �(�3�?c����>��hnlq�E~7D����4Ѻ��,�v�Y�]��SG?!Xpz��Y��C�on+�m� 0�7 e�]���էol�Jx�� �'a��P��Y.<
�Q� �P����Cs�[V���E���-��z-��#�q1�jթ e�fXf��vE��P���&'��+kR.�$H}�el������twoKheR�%���{����U"lC8� �n<ы�T![.A�ku=Y�/�@�X;Bdq6���|��)-6���(�!v�B'�)B.��k.�mW�pf��<�_�q����֗�G� ��Q��T�r�R:A�it�$�-�׆�:��!�����i��U��"7���1}�HgV�U�'���P�����r8i@y��󓚀>�U�Ǆز2cN�p��t��wXi=��\�J7�2�.�6��[�1�>�B#�6�ȣ��!cQ(���ހ��r w�śB.�vV̓"u��_�Tꅝ�&ՏrS���1Y�:�Ƶ�
�F}#�����a�ѕ���y���n�J��5���鲓�ĳ1f�40/���
��p1E_�[DW���1|���V6����O�5*u � ��:���o	�o�8�5c`G�'��y��(�n��.�QVy�"L�<�A���GwQ�!���0���,��/ej�0P8RO$Z/T,w��߰s��o�ѥ{hU�m݈���0V��~>Ƞ�)�\�<U�������7*�)���֥�FSD�x(&����r�"�����v�X3�xƐ�'7����pmY��D��PG� ��e%
�AJ
���f=����3LD�ȷ	|�U�\rk�~�9N*|Tm,;�]�\����.���V�z<&lǇ�m��M�1����Z��j���PH1r�&�3��4y���i� X�θP��}a���ӯ�����W���5Hʿ&+��úN�WM��������a�hnT�=�S���t�%�Dэ�P)��ջ��{-��m��:麅�lX5Iu�]�1���4��p�O)�>���ܻ��&�%����Y�}y|E���MԐ�
R>K�@��I�TE-^�2�@��w+��b��񺍚�z��(�8*4E��#����Tn���J΋�*\ے
~��G����藴�7�0���L�TW�!�>���ԉ��SZ��f0Z���;,�sUH1��:s�mU�{5Cω��{_`�*�O�$�r�t&���ä;_�O|�#5�������	98-��I=�I��BV6�!�X?���Q�Uݔ:���d���e����ےh}�24近lfa��f�ꆁt�;���\�,�=��������o���%6�z��3-S��J�Z�����(�>6�f(5���u�˽�rh���+ �)�@ʓ���+"�}N��
��R��x ��8N�V�PM�=� �I��(�#
o�`ɣkn� ��,sڿ�|������z��L����⌯���?م8���&�l�k�} ��lC�h�!�]���} �h.��n����te��7@�c[����n���Y_���'�9�e2�F�����r*q3������H�߈,�
��[{����)]��#�(��d�:NZ]�[Mzu$�3���8�1�:��ռ����f���V\b����f)�ͅ/�q��_eÀ��'WI���p��@DߤW�x݉��g=��=8u͗�:�,�̚v�y�k����p�- ��L���T��0�0@�10�5�̆�5Ds�e9�5�����4�K�$p�Vh7"�K�:kV�6��;FϚ���V�: �b�M�L�������/,c�����8w��Q��B`#(�E���Wyr*m�(�DQٛd�oKb�����Gh�0�وykJ�\�ao,)��/���f�@W�3��.�n��浾��#DC���=֙��(���L*Ƶ.�G�z��>Q8�W��T��	̀�+��q��Aԍ��7��6�S��?�}����4\I^�p�+%�k'&g�K2Q1���d��� ����Xjm=]f [V�&��Q��c���o 7%��~�������46���	�<�&��9������z��G�hr�3�b�У������J����'��{��d>y�krv�j�q��H�h>bH��ކQz@hH��H�4�M�� �4��?t���ح���E�1��lj�=���mI<��c��W0]�I��:�ݓ�oR��A�e�p���^��bsu�[����;�P/ADں}ig����ɗ���x�ߚ0��g��4���Ie�z�i#�#0�^+X�}����$y5����G���b��j0@\Y�u�pٛ4`��t��-E��)�s�A���<ߺ �eb��ГȑҼ'�$c���a	�m�!a�aVt(���Y��������O���@��YW����6��ų���˷94��/r�w21�3��
����;�nU���V@핚�t}�6~���w���3�؝��敳ʻc�x0@�{�/�!B��$�9��s�-.�[~q}+���r���(�`�VG�k]HMF<T�#��8V�NG-��B����I�T�0�i��w��5�K�>9SE�O�N�Ȕ�q�V։s����]�qBMp��̼��Dí�N��LScr���B�`�k$uu7��\{���#Y ��w�)o�<��q�_��:�zP3��Ҝ���;�%��˜މ�!L��Q�tƄ�T��-^@em<`��ރ��|.���I�|�[�B܅
>q�_UÁ�a�_��:WU�!������!d����vfM|�؁ۣ�_Zz/;|��>v~��(q���ٝ��<w#���*��?���#P�uki�H1t�G��i�>�Bә��!V:��gJ����}<<�����b�sF��?��i����1���rp�$�~�6�Bj�Q��#dO)�܇m%�ªN؅ϧ�lceQ�5��_t�ܢ�ͼ�J���3��l%������wv6�F�*���95:[���$�D8#����g�B4�K���S@�v�}�f\$á����i?�4ڻ;��2������8��&噖3!c���!jP����k~P���fx~m�o�uz��u������T�>��y3�2h˵i����-�Y0�|�
TQ��#�	[�Ϧ��G���B�c�
�]�F,���9tʅ+�L*�W|7K��Qc��d�Kj�ƕf��T*0�|�.Jrc6jN#OԊ�<��	���HO�X���ާ����ja��[�q׷��̀��C�r! D��l4�EV4�|��f&$�\2�*�R#�*̆
K�M�b"�|8���o��՗%%�R��a���d�����|�I.!�͈�B&I���N��}c�C���� ������-;K�ϭ�w�$��*H�}!+O�s߻T�	-s�5E=L�֞�]~l��	���tHI�gۻs��Q�V%Wb�z܍ϖjȖD>���X]c6PmHM y�i��6�w��6�≇8��P rc�B�ֿM��UX�iEv��7
!Ϯ����?f�o@���5;׻��Ts[�їla�ē"�35kO&"��w�ī-�=rZxY�2t� ��l=]���+����P��`�E�����~V��U.�vI�.����j2w9-DL�
w�)�%Q�y������ƃ�<e�}���I�%�3"D��k�^�xZ`7۲� $o �`��H����D=��H���b�z�M�_��>Am>AKt8�хgw/8�9�dC?v�q��\uM1`��k��h��"}��R (��+�l�}Nm;\�c�:_D�9Bĉ�j�>����6��
���`e=F�Ӵ��;���f*qK����}��H�M�t�ì�k�A$#H�5h���o�	0e4hH#pi�D� O �V9�f������K����sa
��\�~o��-������'�{Ro~p̿8g�
kq.���-���O�}�P��ˌ�J�<�A�凱�V|ָ�J������uտ�"��ة��lyS@L�{T��a�T?䩚Z]�l�Ĩ��v<�����B���I��Y��������Z﹘�����T;�&9t����5c�v_p¥~)M�\���J;މ4K@C~I)ظ����#61.S������:�DD�>k��ȃ �����n�X��� ���@�E�jUYQq�9�S�>v#"[��N�w�n#���K�����w�P���Q4[���v�!A:3����3?���^�uMI��Ny��z���-)�����~�؊>�s��g�g�1O�ŀ�Ndo�;�P~1Ԣ��{�m��H�@y)?�yxR:4h�դ�	/l�5dƸ3�BN����#q�HGU/3%-t�yX�h�&�:�H�n$N/5�)��Y�$9���[�mn1+���bN̞ժ�E0��;��`�h;V���{(�/��r}M�|~�<�]X��Z^�!�W�S�Ȍ/1�>v�OSrEw����2\
h$Y~V�`�e>�?W�e�qQQi���v�BAUKL�����$�IY�����vϿ�������oJ6�:�w?!S3�5�a���.���U��r�s�:��
��V�~���!i-m�	�j���,>3݀?��b �Ш�yf�W�w���R>���� $4IL�2�Z�a��x�t��+� �(��1&��� ���z�:[�싞DM����JK��Mo��L��Epü�.���q+��p#���6m�.,߿e^�01�/�Bd���W�7�
@N~��p:�/��h݃@Q� �Bun�@�<�ѳ�B��扼󍚽G�E���> ��^��j���S�;�@ò�x�x�� ��sw�V�P��T��D^�A�_�O������b���)N<A��׿��u�j�1���=B��t�����p��qq����7��%���? �.��ϒ��C��~��1@M:�oB�`��*�_O��Nϝ=Laaϝ�Za&�B�o�:�<��l�l�"��B_'(�����Eix�[(۾�e���z���t�'f��qK��C%�Ы�����zS�Q㏒>#D�zK��ў��65i1+��X"1�w�zKw��D�#�ڦ�g��{��;:]�)V�O�*h4:*^���e�J��i��O=q*"+8Ņv������u��������Q�+�["i)�E���N6^�y=��9.:+C����ZĦS�ڣ�O�*g�˯�2�#��T��h�J!�h]���y�H���dX��k
�R;[�`9/�.@ؖ��,/�f�~�R"R⬚E	�͓���|�/.�K��r��h����'�̢F7�d'ޣL�}5��?��~
�B��ݛ�<c�]
�L�� ���w�%;P;X��>�}�WKh��7-��k\S�E{"<&�HqJ*U�ص��L���6/ݏL"���^��9D����+�*�����ܻOz��t��d.���խu۠S#��7"���4C��I�,&�N|;�<�a�Q3�P#H(�wwicN��.�5X��y�<��: ��玷(%�����l����c۴(J��w��.y�@.N��]'��V�~��S��}�Z�z]����Okgv%�r~��`�7=P���>s�t��\���.Ly��ڡ[.X��7�vw����,����iNN�����2k`-�1�T*�N���?�q�I�P����@'��@��A{���Ѝ�_ZJ����{�u.����ۖ���	s)(ܨ�d����{)M�O��ῠDxa$��Y+��ʕi�ȝfPu���[�\uq�~�D�������'2�E2��,LFn[G�r)�(�o�F�_��6������ꔄ��E��S��3���ޏ7o[�{���!ny�P�o�1U鼘����w=s8���
�N�% �q��|�S��;��Y�6f�ē�{5�eLui@ٻ��r�f�?�77K�d<D�:�K�#��C�^zWC�".%L�<�|ԃ��!�-�i;O9��mR�y���
��]^�E���N���m���J|%��E:�#Uqb7�����ն�e1@ʵ��J�lw���V}e�&���*��"�K�p`�\��W�Ų.�b��4��jek@���:�ٮ׀~�jvφ��������"��1n�kb]I`��W_��5<Xl�g�_��7���ރ3��Yy��p_f��;����n������9�[��/�I�
��{���,��eo֪�F���4�Z�kF������t:Eʃ1=M�ߦv��f+[�>�?�ao�3Y�|�ha��B�����W���4l+Үμ��N�MbO���=��)�r�|�{�A�k������M��p�K�Bv᱅�[VO�ٯ9�(=�g�S,���ԐRC� ?���.� �S�U�����/�I0�'�d:2K��u�`����>w�0��3�������ӗ@�P�XL�#��i�묳}_���}n}�OA:���,a��-^_���n�並��eZ�3�gcT�u�8��y)�m���G��B
D/�Ҏ��U�z �hPR�'�TD���6�,�QO���?�&�b$,�F2����>���a(����_��[������
?�+��(,�8\i01��UeU$��gVr��m�!L�j��M�^�UF�`*�V�SӰa^o�O��9�v{�#ɚyC�\*VA���6���}����&Ŏ��#��%�3s�!Q-�vSW��?�z�+Nu	�������~̈3Տ�m�~����r���d)��d���������g��2����W?�	\�e��?�7p7��5�p?�M羟�;������_�!�2�5���I��=�����RCi�i�ԫ�sa�1��<�$gr��0�� 4�E���*�=xS�-@���#3K&�4Fb���ٕ���A>�����c��j�	nޛL
_��x����J��X ��3�=QJ�`���>��lG:��0�qD�8��*<�4��Σg��.�x��k^tQ�dzgf��E��G��