XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Sl�Ch�ƖK����x|Et�d��F��S��A$~���E���"v,s�0���3�׃��-���.����#�>v'���ʀ���xㇱ�^��{\����jr������wDww����!\��\������_�?�T(J���̜="=O�C�����~
Rw}7�]A�HU�1�9(��Z����ԗ3bQC��J�J�,�ۍ����_@�?y�3�L�j������ڒ�t�N�-h�尒F��Z��q,I�`U�޲�#r���ڣf�,���N��`l�P��*2!�A���BQ4 ���u|��ۗ�q�h�O��}�IeI�d"K�
U�l3�!w�_�����n$0�aKs�}��x.xI3�~��>B2W��M���5d��)��O#J'{�~R=O�'+�j%��#e�um�H��5c�r���㟫%�1�XpPv��-R�y�r�?Vܔ�k�;���������@�[ϙ��#N��Ir
3�@� GG��Y�u<ER0��Z�c���[���ݛc��G,��+�'�nMy����L_�t]���{(�P���T2�N�Ƥ����-I�bFH��@�Y�5��'�X]�%���C��7:�=U�u>�`�1��e���{��
�_���(�MC�
���h�����h��]s	�j/xWF?���w�"j�l�?�{
�F����-�$��nR�6��҅�'������@F*rW��UL�f��d�� H
fz친�0@r�O/�E��]u��^XlxVHYEB    162c     850��%�=1��ǖ�P;tga�'��f���ݕ(�#T45�~�U�ǗE�| !G���g���_Iiy���";�ˣ��Ā[��U&�h��g£��W���lÆ�>���i�g��ĸ�tCis��Qm�C ę+aGB�Q�K�~J)9+�4+��ޣwh��A�aUu��LL|m@#��c��U�
A�!�UM=c��)�5��|,>)���
����$?��x�ʚA�y!�{5փ�/�����m�]���0@쵓)��!u��o��3���UZ�"��h�hznfǞEd��R5so>=�{�)=a?��kn�J�,�C�"zb��������Qj�p[�E�&Mㅍm�j��Z�Ӌbkh�6�~�#�fGb��r�����
J�]^��L|5۫`��ULw��G��1O��^|�?U�ɏ.�����m��C}�Gfo�����+��Cţ�1����Ig�a�?�����tN�֐�H�X��8i�V4���g��hnp��ֽ"�De|6zAqV1� ��S"�&>�3˾w��r��Tߍ�ƒ����L~> �4�3��'����T����bBΙr���Ĥ8[��= �F5�C(�f!��`�� A(�l�~e'r�8���T�jb�q�6,g���9���S�m�F�T�j�)�M@`��S3~�����,�,s��6�Hu�����*������~'����BQ�0�ε<�G����tp�{EД�{hO_k/�z$2=nT�{�r"� ϏT���d��g,^�/�����߭��ԇ��o^�����@�y�!��v��G��Ĩ��
�Bq��ީm�T} F)�B�gc˕�U����(R�\]�~a���\��y2�h3� F(%X6��+5�;�rץ�x�]���!��K����h���q�90�_�yo�sia&���a�c	�ҀJ�m<Y{�f�6[���ޞ�R���m%ݎ��}Ԡ��^�g�����v<�+����k��`TqW��=�C���J[�(��Y�'�|�����b�m�������c`�SG��E,�-�T��3�f	wKc�	��:�jۢ^n~��<��-7�	 v8I�*��׃+��`k�۰)k�z�6�L�R�D6����3J�]��M����CI���^hl� ��Ǐ3��l/�9�,��Ƅd.�%�����c"���B�5'�z�iC�L�$��T�{��(F����~j�%?�r��/&����T"��]$~�<������bվ��`��#� ��[�ڰ��';1aګ�& -H��o��ӏ�'�}�FDJ"x��E���J5%e��$9G.�]u���(k��b��<���mj���ɫ*"Sۺ�/DCw�t|y�;�Ew=�Wu/@�L�1���7��s��E�k�`��4��ͭ��W��\��ʫ?�f6D�ofv ���m��������~jk$���N�o�@@H4���݁KL��I#����H����_|<Zbǵ�ℕ5H�y�h��B�c�4
j�i�'����hOv�Z�)�.6�w������̚�H�%��K�A���&R��A�r�Y=�h��)����H��M�_׾U��pze}{Vہ�����2�B8��FE�*��z�1�dui*���='DZz
��c܀Ӗ���
�W�M>trt�a?2TC1R��PW�]�r��]5��
���BZ��|�c2�W|��`�!������sE��$M}�Y��e�#�:j��hW���ύt��>z����Ξ��3���K�g����rnu�W�ϕ{�QC����ʱ^x`�x��\M6gu���Pei"�;ϓ���;6��]p�����Zyq��{��t���;��$��O��T��*�r#h��x��H�3G}Q2YH}�8I�����C��ę�9,P�X:��-��O��A�F'g�"p h��?5 �ͮ�Nq�uS΀�x�c�9Ŗ�%�A�i?��6���@.�y��ᐖ)"!��uf3V�(³�d̬���rE�1hF�}����_��5���a�i,Q�v�JY��Z�+�x���`�p���
����QI��L�J�W2��<d���o�t��0�2���1�?