XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��yh#=��	,u�S�#!�.7��& b�*��u�}-�\f��YK`����<��ސ�ƙ����ʓ������p��ˆ���3E<A]�W�K[(I���?�w�L+?ou�'����3�\�_��=��A��|�<�C.���`5fO�nOr�F)^M�Ͱ��e�e�TM�S�! To�n)p9��qBTb��3���5�`r��5zx����	G�<V�6��vP��>hѹ�|�^b���p��${�[~M�m�a�A ��d��C$���a�pL{�R��Qc�x�3$�ك�N�k�@�u0��&���t������Pw�<�R�Ȇ@<���ʘ���N���l5�؋%�(�)Ѣaz�i<�Y��d�l*���f�~���9�Y�3�B���Ke4�&^��,������f�σ����<C`o�96��g��H�S�~�G���o��f)�.�ǌ̯��629^WO�S	%���t��������0���L��8e�?���aE��*g'ۘ��ddɛ�&��~��>�	��a!��a���"T�%�z¥�N^���]kP��ɔH7��B��왯�r�d�K�!W�y��z7W�{B�����\�kl��B�봲� 	w<B�����D�ҭ�x�W{�Ho�E+�h4���-$q�{�F24�,M�y�@�-��m'����bHe=�o�j���&���H`�Y��2�J�R���~��.6�0%Z���m2u����eklr6l�gX��>XlxVHYEB    3099     c40�vǶq�g*�Q9���*yP/0���Q�9�&���
�a��R?g}j�Z>"?�/x��?v���+);?r�t���b}��@�u�~�3���<�����ህ�I�����}@-�D�Bi��t�c�1�
ޓ�ޠ�2���ߩ�lt�3���
�~%%Bj_�yL��?]�G��a�ܛ��h�؆~2{�o�rX-@L�8G�>�4#��T����-Ҷ(�ŋ�!r��c1��=�)�/�ӝ:��������v��w
ѡ:e��4s)&��Lr���oa��0l� �~7#��E�MxӿCo"{���&���J��2Dw���H��q�9����a�����i$p?2WJ5fP��xND����L��;�8\��f`�+�$Yw�uظ':�V�lޔp�_[O�� �և����fnƕ��NвI�l�i�s'��[XU��j�x�ױr�b�w|��.`�h�I�2.q�bX�p}D��]�-qd���$Ok�_��7�X��N!��
�>o��w���^�>w� H/�q<�P��6����qJQ���O�K�}Dz���V�l�c���[�{27�~|�y�д��
WXϰgqv�M
���$��7�LDK�5�eWGJx0'A||`�����u���	�q7ẙ/�4�J�A~Q/GV��c�2��`_��$چ;�����|"�|襁���N#�ܩ?�b
>�:�0e;��e���/d�:���������sgm"@������
M+��6�O�m�x	;��Tcҫ�S�2�^��V�]x�V<�.�n�F�R,��w��)��%�D�E���duV��~�dvZ�n�uR�W��U��=W��R��E��[ߑ�@8Cd��v��<W����L��"�@���GL�^|w:?1�@��[H,�*Gz����A�L4����,84�@��}���s��W\��,jO)����W�<moo��
��p^f5���Q�ZQaֈdw�_�.�h�h�Z��>�	i��3/���M6f�1DYD���=�*�@o�o�:�̲z�6XD�רj�w�h�u��Պq�3�2�rm7A8LQz�-�KJ#m�HB��s��t6����-�Y�
������Ӏ�ndѷ˿XBk�	H8�xM�˵��?_9�4������ ]H}՗�+ Y����jM�Z�^\M��dA\x�姞'kW�R�.�I�E��A����2J�̀��e�8���hw]�]�4�(w���"�o��G��+�T�=��G\�����w��TE���r���ZG��'t�Z��o������f�������{�G�0r|����n��#�a��?S��(�#x�vw�	����M��ѕ�8�D�yw���y�Nhڪ:�f-Є�����9I�����gO@�����즷�{x�$�$�������!�X�a��5Ŷ՛�Y��V��v�-{L�d~�Q2�=�����߃F�@��"��7�0���d��͈W����W���H�cz^��:Wt�F|��"�E�����ĳx�B�sԲMmK���̠�"��"[�a���c��y�xoO_��,��0|�#z�m�@� �]�u�3u�� �����D��`��O'F�nQo����$|Ѿ��F��D���b]�CT*2�m�����f���_Hs�S��ak= �t��&Q`8��5G���c��SO����r%�����`>?#�*N��F��-7!�D�w⫖�!�P]�LNePK��s��ɐ�t�2b�u�4����Ϋx�p)��2��,)bf��xt^Vn�bux��b8g�R���2v���I˴ ;��ˀ��	�ݮK��)��?�V�wM�4:�����wQEy�i��Bg��J:,��U����M1���1��2��H$`v�;��# �$�H��v,��)t���Wa��]��c)���ӿ��naJ�.�CG�� ����}�����m4<�A��-�AB�X��ǩ��[�@�@��!!2qJ�OQ oż�z�hUd�;H2����I83�3d��%DizI�%j�4|w0!�����Z�"2��#��6�V���Η�Zշ��v�,�=�e����6pByVkW��*V���J�������lf<ر/��t�c�*���g��՗΅*�{���녮'ib�H��bL�;e8w���0�L�X���;s�y�|��l:����Y��|��(��/ ��[Ċ\�>�0�@kV�uXE�ĩ�����ö �|^l/�2x��1�K�j����2�sW�0��9@��Q�9$��&V 7S�h��iď�k��`$�$��@۠�,�b#���n�Pқ{;��^�������U�� N� �y"`�DW�:��:���!��W�^<�h�����Mz�v~���ഉ����l�o�ڲR7�LM�%#�(�|Aӱ�S���#F�]�J�X�	K\~xyK���[S?#mU�{i!%�X��� b���?��~�-�����g�ڧe����9���jF�gZeL�V��f�/�r�q��������@Y:(�y�zL�@ݓ �J�d�e���JJ[�Ҙ�'�+�F.��f��Ѳ�x�Ƌ�Q�j�0$=�c=�>���aK���ǟ~:ժ��B�xB��+&⯂�0Z�f����7s#b
o-h��L ��@�,���}�𕞾M�^pO�y��I����a����.��k|8�M�]�d����g��W��/�օ�e��o����v.�����}r��Q�Hs#ň[�om�*�l7��ڈ��n���IT��G�5�B*���	�12y��ձmWy�%����	!�����.-�4i��Oҗ)�����Gf��]7R*����*�� ܋��K=�l�".�M����&�#�"���)'��ɹ c`�ҳ[,-����C]9�#��s�I��D�%��E�� ,�v���J���ŝP缽gF��+�a���@Z3��=p�(�G�B"��Y ����C�B�bG	~����$��`��O�-��Y����h��1���Fr3����
�U��"T��L,�a�ݦ7��<�D��v=x�ɥ��\n`'/qڪ)�����Z�}��E��[� �zF]ݢ5�K�����7�	�囱t~ög��f�;