XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E�k�c��n)��4 m��.<�2��ܲ��E	g-�.k���#?=\�/�G��Z�~u�0��=OD�X.&C6��m
!���谁s��8F�hzA�617!	t�H(&����}z�NR?7R�EwJ�~�0j�=�qh\>��yc'�KG����Iq��Ms�C��j�KbI}u�<��xnP�y�n�>�m7�8o��֋���	���bz�&︖�.��d�%H&̠;���*����x�{��Ӭ�;�Y����ڴV���h 0���+�EN���vI��]��p	��liZ�� ��w��L���ɂh ��8ؾ�k�S]�5y�DH��_T���r����hB{�ugI��
.�3���+������G9��"��$��:[��	[*�Xp��/u(/�5��6@��#A0��L���(v�m[�P��f�J��-�R���/P��TK���u9����\2f�[��ͫ���`��ѮZ`��e�>2�~B�Sq�`Ư���jv��{j2t�?^�W�Km����{w�upM����rx�Y�˺�g�A�IR��wN��[�إP��o��`"�?*{�M^����.p_	�Z��}F�M��;�=S�=��Y%�Q$����a� 4{	�������Gm�x+>a�B�ߎ
���c�_�Q~���4B4+�d�1C��`c�n=��ԫ��#�7���L�!�c���,\�����޲֠s-������\��IV�oҪ;ؒ���CK�|�XlxVHYEB    29da     af0�3��I��ap|Ka���Y�glR����Ek�j�M�0��3<�DY,&/Pye���a�b�З��Q�ݰ��M[�vo��Le1ã����⻋����EZ����$�ޜ{m
r~bxi�:T����zfx<�3=�=.��Z�ރh�7�$��<t�
&I�h>1)/6c7��k�U�����՘h�{�����I�/��im���WN�!�;�������������I����0��~���"G�fm����x��Yo*#�PɲU��E^v�ޭ�ｋ\O����ݹ4f�k-V��3��Qn>�[�#_H%�������tK��������f�8�;���5�	�`������١�J���%U�/aQϛJ6`�R��4�ȥ`� �Lụ��bo&��)tnӾ%�2Z�֤0K����u������`�k�R�5KĴU���%��]K�v�,~�Shg:�H޵�R�IL4�Q���@H�t�t-?e����,��
0�~i��r�W�4�>%��X
����&[��!��c�C��+|�������  (]�M��{����պ�¶Z�xrfd2�r]��Q��:	�ʂ$��D"��$3rD�𙼥�4�KO���Wt�����=�����$�*Qq�㴓��e˓yc&����!I[kv7�M���,Tv�Y^���W�!�^6� Y�~Z�����Wlx"�Rܧ��.���(�G�:Ϲ�����[Ʃ�ܡ띺���D�بX;ӦêT�2��8�/���t��7�z��;���0��O�ۢ�Y~XGF6`Ik�p߫����W�p����%��?Z��؛H4y[tb�#kB�n������,����̻���C���LE34�q�H��ޗğI'J�l��*��{��_��$����o��iGK�D���f1�nG�-��P3f��~H��u�쇣�6\��"�<�j�]X8��<�t��+�r�rM�fRм��ž��T�b%�ί"g0�O}v��Z�m�cϿ����XL�.���Rqb���̖���ۣ7��\h�ɫh%��^�o��qK�S���%nN|�O�t���T�i"1���4AW�����5��P(�8����;Cs�_�.�K�G��U�{<1,ʻMچ�#���-�ǚ�K��{��_�����{��!�HfQ��}ڤ��c�yl*���W��WyH�3�D��!�\Rh����^�Dg�{gÌ���sK۹M��)��&��L��b�^`�]0�=��AY���J��:�Q�Jy�Dv)�
��/g�b=;A��F��4�Y�1�q`;IE�}\A�w>��p%y�P�������{}4�E�.�#�$䶠�u�	!��JN����;&�x�� �tT<�]b;�H�C�-��. ���rh�0qa�}����JoQe�.�`ȝ�.�>�a߫��E��,�@ש�����@��WOM�5q���1n�� �1�²�� JY���A�,i���}��Q�P�m����R~p��ı3��w���[��PM���Gm�.��{H��=2�
�;ެ����e��H���2N�A��<�2������ʡ�"YM
*�/o�u�Z�<vJ�Ŗ��`��[L���
z�,俈�aOˬʺ�P���!"�m<�S�f����/�����UE���^'c� �P-|iwu����̼(<$�(�dJ�p�L	����o�zB�HQG�6�W׈#�~��r��ERa��ǺY���?�|�AN�u�A�`ҮN���� |]C8�9A2�d<�K��0ŉ�%�6�&4������:���E��{�2�Cl��#�A��Y��;�YBX]]]b0�|�^����."fb��~a�q�5~9'�X�u		��bQ��tt��?��t'�V��C��;>)T�s�hjr�N
��yp�es��n�w-/��`��>�@�&�މ�|&�PH�]:���a���ʉ�O؂  �6��I�q�����1��'?^�w�/yi�|?o4���0f�}���&�Ɍ�?����P�p�����v�b柼]K�oy6�U������Rؽr'XoX��&Cّ{3 �����w�<mi>�S��ڂQ
�!8��0�����uQJ%�G����	^��2��|eL���u��:��j�����iݣ�Lu�Θ0<�;�b�a�-L:���G�^kJʯJ}�h���HLڪ����a��V��|O��pD?�{{�7ҝY�!���d��ڔ�|���`��| m�#��E��S�W���=ޫ�Ӆ��'��<&�؍'����#o����|�W����D|qk�k���l�<�3���jɞch�l$�8@�5�XvE�U��}<O@�ƺ�M�-0�驣�갍Y"_�7��#�"�;�N��7qc�2��ׄ*��?�L��ڽ����0Te�}A����o9�6|J�mf̴��ϷS!b�W*|')�X( �Ѡ�V�A e�޹��X����".І�[U\���2���g}d�F��z��_��]C����ބ�Sث���
|������;�}�Lh�Y)�,�3,�(�0J�w���C�[�4�b�9���2u�F��.x�:�Q�oHG*����\N/5�1�@�n�����M?V���U}C���7)�����?p��)�<��13�̘�>�#Oc9K�k},�-�Z��gN��<�������ۇ��׏�����w�rjm��4�1x�Y*pp���h��2N��r���-��WA~