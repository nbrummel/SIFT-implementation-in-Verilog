XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���<S�[��c��v7$����K�׏��V+bZ�hGG��k�ց�'��ɡҋ�b� ��J��yC�ܘ@|��W�ۘ���H��|:�]b!*0�)����P_@���"��}��Qo�����hM{����Л�������sE��4�z0�jt%R!1�2k�z`�~fk����'W�u%���,ٶg��u�o\���Z���^Q��� /Q�!��{��糩�������ߴ#ZA*@���3&����#A+�)�f��^Q����w��0�E����@�y�E�ԢE)�:Y�ݬ^��D���
$���cK���wft0>&��)$IȆ����d��Y����J5^��q"�o����MKPs�����5)BM��0:��m�&������,{�p@�������&�fĵ:�Gi���2�˹1�M��ܖ`�5]GB�0���\d�&�r� �%-\2�A(��^bu9
הu�0Zu�����|P7O+s�	�� ��l@#�˜(�6u|��ެ���k"�TrBtXā�J�D<	̛_�2>)��hy-�Q���C�a����y����%w6d9�ݦz@���=��N�y��ϼ3�ß�@C~f���uD�~����(��K����a����w|� �R7QVy(���r�d�E� ln��;��������h�1�MD��OzH��ô���+3��ϩF(����CWD�1��#}D+fz(��zQGPl=#�uN��#�Cb^��õ�2	s6"N��Cs��:���)�:sXlxVHYEB    1a5b     890W��?�EL�/���;Mh}_$؝�z�[��1�X��x��NLp��y�N�.�@�mh��e���1g��Qd��Z�`z�{WV��M��+�z�L��VNO�׬
�������w����3��n\���'�w?U�,�9�]�:��l1���Nn6��鞛
��!�y�hoF��y��t�L �_�N
��)����B�J�q�9���=o��^>F&�Ė�*?BJ9��g�w�*�R��x9�kɲ��\��Edc>˵OM9��5)�g7�"��ܝW7ױ#: ˓��6"��K����z�b�N���/����ݞ-��	�rG;Ԝ����q���7���ٙ��!��R�	��_��y�Z5ez��f�r�@τ�Ld8̳�+AP"���!��c�T���XB_D���u�޼�0@+]δ,��϶�Bq�sퟣ�l(���!�9�^t�C��*n*�P��~��Sr7IɌ��Js�^Q��"�:yL�e�J��؋dΡ�j�z��%���GolЌ��IBe�eV��h�Ⱥ�؂�t$Ң��������<�nt:;W�Fƒ�z5�g�|�ЍP�mMݘ?N���8[�P0�����Ǡ'��{y��8�D��#�7W�x�[��wG8�������P�@㐁T��JO�_:�6mJ!��6 �-Pe�g��`�hxZ���v�
�a�L�6S�zD�&v8��\�S@�Fhk�<�����'��,�9�E���m.�sv�H����D����]ҋNV�2���(qY8�R������i��M��,���3Zb	�i��?�
x~#���	�S��%g\�@���m�$�T�U�Zw�r�6r��?�ǺC�)����{��~劤��7��$����2��D��a�s�UFD.�;��ן�xלx�@�^0�fΰ�&�G�C�R��S��)��4o�ʯ����^��! ���āS��k@��
+��6!���z�t$�9������%w�_�D�CFZ�D�V��%4xO����#��8T��c4ǘ���bR�v)�ZHo��u���R�_��� �{�Z�Q�=p_xz�� NF��7y��j�ۍ�Ь�K����(Nb疪k��Ha������.EC��]n��u���p��6&��]a'y�~2XKn�d�B3f�ănb��{��j�X�Ë�\yi�X5��Tx^Fm����^�9�3�����s�  �|^
ŒaCNd@4#�{��p��8��X#��&L����P��ji<T.籏��}T9�ȅx׎��Ͻu�k����y��! ުƭ���|4V�N��i���
��'P�{� �)�/�x���1��/��"�'Uzd�Gq!����)i�ܹ���%�q���i����H����Ă@4\&	:�Ń�Mُ�w�+E�Up�sO��k!�*�t��_o�c����޳�)m�u�=�8k٥
$���R��O��4u��>O_ut��h�6'RB	�0�aߠ-1�z��aZ��٥�}��Ȁ<�Ṃ]3Y�S����4�
l�̂jt��AL�S�c�V;s�V�<�� ԚObU�in����z�w*<�`�;!�ʊm�:'+8�m�'���H�|9�\\d�+$>�dsA]���a^�d���={�<I����]U�Ly��6�<H2L��`�e˾�F��ڛ��?E^D�*J6���WP�q��
�?�u�I}���P�
�ݔ*��:�Yya��$�4�ܮB����X/[�>^������-b�����걘�o{?N�l0~�xlL��SAv��á�i�?*¥���g�b�0���T�U�ZI	5�w�}���7G��\�|)�����̵�@R{�-����1���	�a�zF�|��Ă{���5g��n�춞v����)�?�՜s)d}W�PPڊ�6�78����sQ�;Wۢ��F�	�7�q��gŻ��oD0J�#�3^��@�}Pt��2�������^�İB|]]r�_*��Y�N��.}ؗi80˲n-�e ?����_����vo���2Kx75ñ����j���T�<LXgz#n)Q|�&���kw����G-�Z��Q_*�%(���{���Z��R�0@A�u{��o�|��K�vo0�XQ���	.1��-N4is���u�D�ֵ<��&]5���3��˪