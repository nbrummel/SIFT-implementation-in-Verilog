XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��bg�RY&�'��Ǐ�v��r	�?��
(��7s�I�ʿ�S��(�-(����NSt��;$	���^�Ģ�ik�m��Q����ȟ���Wr�>��{�]���VZA
(�N��R�%��S��",��g�Vd{
�2�YSY��y�S�$3i�3�Sy]98b�s��iw�T&�*�㏟��w�K=�C�d�[>���*P�W��Ɍ�&���J>Z�N���[�m�aC5f}LTf�r5Pw��@l��z�a����|��������= aR�N�:a�/��N�B�I@����8d�1��Ab��k�J��a@�U��=c�o�; ���Rwr��W)q���탇��=�s��4��5c`�0Òoe#�Z����e����3��Β���k>�>��Np~ ?c>�ߐ������i�����!�QV)��yD�jx_Vek�`��w`�틷���ک��,f�����7̈TW��6A��u�;wkh�5 h�Mf�4����k�	� z�l-߭b�D�~(�Up>4�s�`��3�Ftt����u���L�Rfv#b�K+oAhJt_����H��@���WI��
 1M���O�E�
 6Ǣ�߈o���`�Q�ǡ���8&U�t�,}ض���^t�7_���jʒ�!!�%G��bY����L��ǘ����X\e0������9����W�� ��f)�Xr2.=��K�eҙ_�g�����#��'����%���04��\����,�M
���y ÝC�Qᙤ)[1XlxVHYEB    fa00    2480�u1Zd� )�oZ�:mbf�nӦ�BQ�$��\c�"����~,����"J��; ��ۗ��cI��'|�U�ܿ��������z�7N���^�dU�h�z���5|߷�aHVB m�&�
F��Dn����cYZ���G�Q�,>p�۠Ԇ�+B��_JI��R��?L�	"����+�'(�~�Zu��(ۜ��+�vlzLa\��`������	��,}X�d�t �Hf�wX�r�'�4���Ol����}��c;��]v4 � 5���C|cyJ�)ݲ��&M��X@=4���#t'*vz�W���X�ɝ5�Ou$�ˆha{����"
�Ц�#��C5jF�W`M'�It8�wGA�"L+ʛ�̚��;��w�e4+F�W;��Tj���n �n�����vTZ����1���ڑ���C��A������+H��ͧ���$#Tb��߫]�m���R�e��dwAS�a[����q�����|�v:h6�vA�J�
�U�$�M�,� ���c��M��Ǔ��cx�n�Z��_�XSەB�(_2�� �p���i��B"�n�H0��qs�
��9�����Ke�HW�����C5Rp�v3�d�����u�����H�OyZ�����'��yQ�XN��ɩ[\�	���ツSj���Ak1]Z�/7�:މ���Dr8�쁰��A�n�� I�
\�a=-�4��R^zl��F��c��<-�0���~�n�K�F ����]N!�\Rm���%�J��y#C�.�9�m81��d�Xh��(�Ώ��rlNٺQ�u��h�Qj`~��� Kj�;��KQ�޽ ���w�k �P9�����ϣ�����;�KuP{�۰�u!N���0�AyKsUk�0_Ԇ��8"ʺ����-�:��hc�S����@k�X����ݢ�$r���o̚	S����c�[ƀ�C�^9��X����.E5�Ae��)�KN܌$�G��#�����#Ay!�#+?ۈC������� �9��&涛��nZ�k	��<;E�x<A�h<�4�O=�D���� �~I�>�O<��n�J6�B.��b�'ݞ��<OET�"�k�ͷ���Tz�lٙՍo^�n��}�r������ߵ��N�i��ZF�&|�nX��ĕ[4�����w}JF$�Z���NF^�H����9�����rܶ��{.�h��j
T�<j����b�Y�_�m��ӺV!��+VRwK|ǝ���4Ұ��n�,��ħ>`h4
1��.�L��E��Kd�y���gE�ƫO�/l���\�`�~��-}x�вV����"?�]2��X���*Q�76(�grYޱ�xZ���U&i`�Z�n[�Q�*-����
Ⱦg-��,Ĩ;}T��4g�����6��u��*1k_���+'@V#��򲱎@Ԙ��o���}���h��o���`���d���X�y�Wj�a[����W��xuT����[��8f����n��<��v�T����,�� V��",�D�����>ԑ�v�;��R����3�,j"ˮ�,���ۍ�N2ڷwp͂Y�}r�A����(_׎xd �qG���IC�O LԈ�ۨ�����:�|�Kl�'���j�{3D�N_�~�{Rt)^�@'o�l�G�|c�Di۴\Ӌ�}�;Vw��%gU��r ��~�d�5WrJ�˪[٥���l��T'���d:�6MsI �	�;�hi��.:����}��Α)���:UW%���i���"T�Y�^I�M��S�����5��L(��E���@�{_[l���,dW�z��r��qq8�D|	�KqAc�2{>�m �KX�Wj0��p��͐�{��"0�nE8|P��Ϙ�%QN���m�9��q�3-~���Q �*�b��Eܒ�dH�\����.�k��e���y��W}��k�ͧ��'����th�D�@.�u7�bX^�k=浄L@9�w� �~q���l֓C����-<}-yD���s�.;���s;Hb3�����h�ć��o��7���{S.��/Q;&�On��{V�����t�n�);��P�g��d"3�I���^/^��1lY*�ot���ȦRVl�tH�TK�k��P�;裼tp�*�*��)\�BV1��Y_��jp�h���H��P���
������Oc,a�DN�[�n1]�����������%�������9���3�LlJ����x�^} ;��	#�U��5�h-���j%��(����mhr5�$P�"6��@`��]y�8�)OV�cŅ�{������w�,/B�ʔ@g'�Bg��d��m0[���5��(��^��S�gD��\]g^�q$a�J�"���Oa{��-�52_�W���YO��a��~<����Zlf�>Bp1�����=���8zh�%�=ܳ $���2�l��Ңȡ��4c{t���R���(/�rq���)=��aW��/�>��S]���l�A(7�4V�Ѳ�qp3�$"3���}�/TCi�*3��`�'N�Ɖ�~����ZhJ<'����6��V ���̺����X��<���V�<���0 �H�,"��x�6�M%��VҸ�Bql�|"�]ؠ\/�1�����ОX���Җg���@̼,8��5iSʈ����V���y3��Jɩ��O��ئ�r?J��\Cwy�N�y�4�u�4�iUq	���TJT�����-���@�2�|�^Fhy��DZ,���;Cn����30!0�]�7����7S��FL�YY�.���sOelX/pO�Mڛ���i�P�x	�w��1o����u�)�-�U<�,V[����X�Ĥ���^�ʸ<���<ޟ]�?I�2r��!Aا1(:��6��7�5�nb���D��m�i������'�<U��`ΔY�0��Id����9���84'=�����Y5DT#�c�qf�@ꄢ���e���+>\1j]c��X�g+y�ڸ|� �R5�c3@�Ԣ�FDY+9����-���U�S����A=P����T>8�4�U�'����K\�έ�Us���@�H +a������t>��w�_�d�ǖ��3������5-�:����E9�`� ���`ӓ�>�r���?�W��:�"r`�a�=��b_,���+>2A� �?�MB~�r`�*�;8r-����i���|��诉�⟉2���8WT&���X���J$1���\��xX�������P���|�O�]_��R�Svv<c�,A��z�?��F��9����4Ҏ��^��;��ZZ 2/e1��Pp��JR�ˌ����"3Q��8��C��]�P����w�*о�JՃB�K^�)`l�rW�h����hj���E(7\D�``�Z:�J�ў��FԹ�*��˚�hԿ��T9���� �9~h���/���_�ƐP�A��j���#�|��kF��h�&�c���ԛ������ Ү�<��͊#�h�ҍ8_g{�J��ꀑ�yUoQX扥�0.M�/���d�m'4<-���.\)�!���R���Č�tä7��(>�eW�����g�V�������3�Jb+�Ê����h��v�5�N���H2�!���8 Y��>�f����Y-�_��;�d�F'b�lu+%ѽ�/����c��~/o�Lrn��FS`��ǒ)d�>���Z0��:�7��_l�G�.�h���+
=�0E�,Ǣ�ł�_vQ���=��Ӵv�4���6Q&�!���\bgOc�!@B;|gI�]�U{{�S�!�9��<Հ)��̎���l�eb�(g3��#�lG�iD;��D���[��B�
v��U�\�2.�m������4���>[�5kE9X��Y�J@��� '�_�s�L�1�(Z.%j}�JU�<���t /�8\��ÄĢ7 z����+=�j"����nL 1N|-���,��d?�w('�h��Q�o�*:��-�@�..F|\�]��K����y���i��Q�k\�C%=�Qca-�g7 �F9�ypC���f��&}��CuA��,4݂�nS� ��	�lR��W�=l�������%�CA��w�
>̔jS#Z��%ؠ%<&����7�[�RYտmN:ց��ã+��Ie��e���m
鮜mpJd���7=!��H�m�o4��l6w��N�@���5�[!�����_�M0o��r:���Q^���d�� z��X��6w�`�e�n���v2��� b�NA�Rg��D��z���aDc_|�<�<�ZZ���������n�D�o�P�G��i��� Q���d,����,��!r{�Bڥ|i*���o\�=���;��5��<6`����'�˗` �����[T��,�X
�2���1gDai�0�_�!���Z�U����y�^�W�g�{�1)��p/O��xu=>���/ظ�]Z{�����1������M��>><��՚zj�4�M}]���x��k���3�ˁ'���*,�qƓ^H������Mg
Z[nDj	:~���s�f�^01�S��.��dj�D��)�S%�S��� ���S�	�P�p��{��@��7���[�_fx$��C$�\�pEn}���q.���sɂF3��P��Q^���#(���8S}:�e����Y���&W�u�(�|��Q�����Ɖ>��*3S��6Lj+"�EuH��|:���1���ܖIn�>ӑ�&;�M+��QF5� �`��t�=������L���J���ꯡDC��=ҝ��;.9�����7|u&žS��K ɦh�{ێ������8L�$Wu�ށ��SlnĔ��������J�X����Q�X�U��5�\ҘO�A���l��k�h�5�X�T�)��U�|	U|�N3�� OJ���4�L���Pxm\8ߙ��� z�� �Uu�䳿*�-E��A��5	��G��=�Ml������瀞B/j �a��U�M;(�o";��qʕ����أ�j�$hW�!�s�:U.��2�@�#y�Y�[#)An�"Iw��*���j�h��>/�=�#Л��"��� �Ӯ�_N�� ��cp��Á>�
���s�v�����Չ%��-6j]�w��]Vz

ɿD�櫼���T�����F�~����нk@�kX����dW��8�7JÆ?R�U�$0�����������}�H�?,�	:S�L"�����m&���$9l%3/ ����/�dw��t���2d!�@��ZQi��Çw�	��.�o3��2h�˹r�����F�e���5��4Z���� O�\�\aC:�[9=;R줞��{qF
�R1�b ���J���l�T������я��@D(�|�3&�#C�x���]�^*թ�X��yJz��u��ֽV�D�ոh,U.��@$<�r�n�ԫO�n�i�踧�]k<.��޿	�����|�Ma�+3a�6u*bb�n�����,x�ˋ�������Z4w�2�fP���������\/WdG�����o ��Z�A|^7�&�t�Zui���o�C2@Y��g���av:b�E�/Z�'F����W��h�9qB&t��2A��J��Mʽ@�w�f��,�q%�v���T�R�?�3���Zǈ#�wp�<;:q���+Մ,�D"ϧPȍO�!e�L�;�̓��K���C�~b�-��׭�x�`�	��`1�fx��sw@����V���j*�f����hDN����9�wR�V���g�
tS�A�T[�.�g)׳b$J�[���4䛃�.zna�j�"X��9�w��������94_�Pb�h���U]����(�hG��U!�.�z����7Y��Z����T��#���BM-�
�}C�z�7ߏ�fVIY���yH�p��Q|p�'�A��]�)}���7亷P��:{��������M�J�f'g�ur5�o�w�1��\(�u��#K��.��n�I��9�/�K�Ɔ�>���a�ɀA"�LTe�d��a����]�jw뢍0�IKZ)�U2�ac��Q֙�fR�����ҹ�-;�hB�/<<�{kS]�w�ş��A;�!��G_�Ұ���r�)��|r%}߱�D^�E�=�h"\�?�pkk;���k.��->��L�EqD�\:6��Wx�7�F�bڵ��J�P%l�m��<.���*�@��g�g#��3'��+��=��`G&�|�?LC����	g���M�G�qoFΚ#j,�+�l��Z Ē�=hBZ�݉�|�Sϙ���c��0T�ȏ�$�m>!g|@�79UM�g����#�d�� ����!���
��)@���VGƐ�T�w}��\�*9]0�{���C�b��~lΣe$(ys�<�]�r?�}����� ������I�6�,�n#�#+ٲz>3�����<;��]!�c#K�|~$7Aѭ��2�S�p��ؠ�������yI�mX6L���7�$;�bܬ�8�I�B�o�v�cN�u�7;#1�`5�0���I�C��K���zI6��4�E����,��}��b�0�Ѫrw>C#&^�\��Y��MGM*�%���i�W���L2�E#�]��Zr��ꐉ��V�v��=;�?C�nM�Aϓ/`���`c�U�5D=�w˓?���m7鹡�mM���f�J��<e��4� ����}v7��@��f/�t�~aR���م���Hi<�i�1�I���׵�Pr�G�W���ԙС���%X6��Da�ο'&�x 1�o����@R�|cp&���׳�#�v�bG_�٭�Q"��?�(�2!bv��5*I�����&���n9$��r�$&#;�|  S�D6�4����ag��cY��Oec&+�]�;���5(����ױ�k��� 赎��,C7T��C�>H��� �-��=MiP7D���ی���^A:����Uk��2+�{��ф�}P0Nr~6�D�Ӷ�����dY��Ļ���ё(9�R��@�4s�{�S'��̗I����"}����מ����7>Z��w|ǽ>'����hiD�&��Y<C����x���H�t��ѐ���"��s�6���ݵ�=~����QM�8(���E%'Nq�^\�������G�� �=����L��zO�[ɔ�\D5�Qb
\���*��y�."��d�\=Ŷ��+���4��z�=�L8��H.qc�	c�D�|�x��. B�Gٵ�Zi��'0�W6|�0~�r�z+������f,�[,Ғ#;�n/��9�F� ��t/�����⣄>����~��T�AY���G�������AK��w�+T����GC��K9vʟ��
ؚ��!G�Ϸ��ǖ	�N��{�L�"d2�o��J'�Щ�b�Tu�#0�w��-I�=)l��gA~�x?9K/Iap�>��i��c�'������%��u�K�k�X�SG�ޥ�+f4`���tn�o���&�v}"�������{+�y! ���`�P�%��v��V>U)��Q���������k�{��QY������Ո��C���.ɬ�/'ֳ4&����d��V)�)l�b���i呫u�u�Ӓ��*����C(H�h��r��Ո)_W6��7w��z}�*��t����D�(�C �R^�D�öxA\Eޙ,x�_.�%�F0yR����kB�sf��L �)7�����77����ъ�Ҿ1A���(��w֕`�W�. ��?U�+��L�A?����g���6��(���$���nn��$��Tl�_k���#������u#]�<�z��q�ej��Og9,���z�?�#��U�0��;�i���d����mM�C�c��o_yLIo��̶���QK�ӏo��b����+
��o^�݀�-����5�Ip��PWV+��o�
�S�0Q���5�:`�z-�U*�c���d�ӗ	�ӓm�H�R�i��s	e �-��5�1n�TƖ���b�	��z�3�]�i���{�X�������̧����.�R�s��$\���:Q^�3�(yA��.0(Ȍi���Ӎ�a�L�ec,�G�1�١y�|Ǭ�D�g�uD��d1��(�Ħ�9�ci��L�w��G��H;��n�t2Ĳ� ֔e�)�Tˣ�H��č�wź�.I��Ҭ�9]����z3�C���;�hH�9O���Ʒ �B�?R���K�ٌz����E(��<�)�Xh�Z��`�hu�!�+kP�ogZ�3,�������[wxaFzcw*�}׫���[N�#?H�ֆ��Oh��+�8�>_aY��@�f�f.At[��p�g����t�_�X-�Y��&Y�1�������9L[^̡����j��Vx��{Fڹd�=��c���;�������>U ���ˑR%�N�+��	���-��ak3�D��!�P�V�hS����4Zlۋ�$$�GS��"(��� ��O����s�)+�ck�K��߿�M�x-I,n}W�L��!����������jd�ˁƆƼ�L�4�*��}]����ɻ��a{��n~ȓ�/�(#[t�,��GkJ�����ph�S���2�Pӫ�'~t�u�C먈p�Y��U�F^��#�S<���h3��y�v��YҘ�(x��n*\���W��,�K���y��+
�r�p����i>~;�Y�Ǎ����O�U�Nn�6�wU���9�SJJdn��ء�(H��m���|9�HS�g���P�U\2�	�&��I����sr��de�Lܹ���h%�����M�P���LoCf4��� V�v�	�x�5>(�54.��c^��t���k��@�����l�v\����q�mt��d.�ʬ1t��9M^6�Q�Dy�\��� *���46��;�R3��N��_+��<�����@R�>�C�L�l�J�Os��Ÿ�e���'��e����#A\PM=�_Í�U��z}��T��A�^@��n���,�DU�"�� *�>;��X/��U�1�T�cK��W= �G7�m��F�ǰ �pʄO�%1`ρ�@.�Y��>X���f	!��,�^��v��/��c�l�CxzVT̝v�� ]^F=�O�&��G����Rێ h��KO�h}\�\�� �O`QEڤ	�wݺP����#+�8�-CT��<�E��h~�l��ʒ��M��n������`���d�&��9���R�M8J�j«�: �n�q=XlxVHYEB    964e    1150�s|?5nKK���P4V�@���{�.���;�mѨG�&n���Ǩ!���4������N��"��"���6���:�XEA%�H1��bVt
�˷��4Xt��1z�6�����W?��?�ڗ�4�3���2�u˙��1<0s��V����*dr܉�Y@���D��ſ�1���Ղ�ⶔ�=i밁s��T�q.�7Y�mF~􃄼 ?�����I���B��������]�]��.�h>�^��%��``'��ۢ	���ui{5 ���!}�TNH&�Q�X�ju�m�XD�+����&�9�}�\Ѻ'XgZ�t���/&�2o'�*���)�0`�E)C"4P�B� /�����f�<5%�\�k�eQb)8/��GNr��R��(RD'n9̋��c9Z9�S���dq4'�7_�yōR��C\Y��Y�8�3��T����\�ě�#)�ѷN=�~c������e�w�$��U甁En���{�cFBk�j/W���P ,�0�Q�v�|��ɒ�~?[���V:z��o2����PV����
7~��@���t�{�f��n�Hup�'� /��Z\�C�z0�-���Pι��	��7ʍbG��`!�� H&���3Q)v�e�`L���I���w�̥�D"�9m�6���|��PRoGY ���q�:�V�T���6\����b�36[��c��XG�F�>�o��SA
-�n�1���?�g�����8Z�E
��Xr�?�?����8� W��N��S�H� Y#��� jnx�ƾ�[�P��Q�&/�l;��H��jJ��8�&�2���!�n�s^g����w�#v:uZ3-�iT4XO�2��؍C�v&?�~ �iNص����!y]�����m����_
��������p ���FL3O�ՠ�;�����#.T���[��qZ����%�(�]g;$�v�W7��_���e�B��3zܟ�2/΍���6���JM�?�`��:�$O��٬x�t<VrQ��*�M��R%�	יj�n\�D5���*W5L����Kz"�w�(�&;}��=�*Z~�{������Y�7S��*+��חiOuR�v�v,z���t�h�=#�'-rx��Pw��=���FZ�S���ǂ��t�ۣ�6�Z<ڸ:g�b^�w�����-F��5�E��'��S6bnrPFK�誮^��{����4�ql~���$X@&��,��`��ŷ,J��� ��'Ձ:�NW����J
��b�Σ������q/�F���A�S����v	+Gp�o���jWU(���T~혟���N��-�_.˯�Z�i����L5|�<�w�8��Z�z�:)j�vI6���M^/V#�?r�_Ӛ ����ư�-H矢_H!6����|��>J�����J�l�� ��J�(w�(|p��~e����vj��oץ��C�ޮ5���#��yIF�*���U���^Y�>|iJ���o�A,�
mF����6P��z<%j�<E��J)�bA6%L�7�FQ
>fl^�R��L������^r�iX�1^�*!^��s�?ˑ��-��'�̇�B�+&�c>�c*��+U�^Yԫ>-����r
���� )'�_\Y1dY<���1��`J��ik�P��D&xY���ޫ'��L�]	�);��֘ef������ZW��P]W�=N�V~�	
��̀@����p��"8�K�'&	aL�rH�z_� ))�P�SAzt6�6�a:(���l�΋�����7��2�/�}\��r�)��:��Q�{�]+K��$I*�����HQ�0��_�K�����Iu�Pr'��ਔ9��d���V]������j���`~�G�x��(=0_m��GC̀(�<9r���{~-
�*�A�o;>�/�rX��s�-�r�GT���T��zς�*,!A������t�Ƽ�Z�����-zR٧��:D��K4�5�m���a�Y=5p�5O.���K9�c�u�+�u<],^�TtG'�q�w< 
J��<yK/�J�� !�8�*^�岴��c(�$.N����%���5?�CD OH~|+N��H���|��UF��0i��Z؆�� P�+���8p�ns=�l;�e��T��n6D:�h��Ld���$�}��[9�GsM��?�7��R7�-��I�����i��tSj-s�N�\���E��A;с�Z
p���&�F��]K��nK;]0�z��II�� �.K���j~�&o�K,t/��B���4	&b�U��|�o]G�>��~�� �l�Ñkҋv��\��@X1Gh5n��)]& n��ٗ�-���P5�:{�n���o��\'�Qd���U�L���!��e�4��զ#�^�v�r�l1�����3��!K�-��u8��l�6kɭ�Y�˘-Q��p>�����[Eӷ;��R��v�����w8�f��;k���t)��F�.��Ƣ*2�Y7FŅ�� =-'�h-̇� f�)($�;~RMf���&�b�&�N����-���&�]�sk��3��E��L����}��(�Xˣd����nT�����$//7+�ۂa����.�/��k6X�?�J�Y7��pd������"�>$4ggw����̱���w�Qm�g'U����6�H�s��6%CWl	B��[D|͢;E/��ʪn)7$����,9��A+,��,��̂��QS��%���жnXO���Jm��R���o�r���o��|���+�=�0��؜'9H�ۃ����O�yE��&6�<ꆚɳ�+�;�=K�=�A��])x���;�\��O�2 )XF�����Z}P�B��`��᳈sAn�aw��z�x[�V2NQH{XoO���B�c�-X?�w����i����QTr��E�i��(F�.�rja��-U�.pf��jЋ�����cL���s�`����jL'����c%OYG�8>⤇�b��ӣ�.��"�X�9�����f69���'��� unR�I*��eT�OP%��4�0C���ڊ�������⨋Q���V۟�h9��-ZK)��ol6}T�"�u�PdL1~�/�����dg��ԗa���y����~�f�����X�%������vX�d���$�A�Q���Fs^xb
!`�=Q��T>�,�$G��N��8y��3��pVu���KF[ף�����Y����8&o�B���L��gAoo���HtSd;\����@��7���'$Z��;�W��JxP���Κ�ϴ�)��ڋK'ڐ7�Z���ږ��)oJ��a7y�jD}�F
n�@A��s5Df�Gq�)�B[=n?u�#� [�!���~�gV,��vl�����zW �]����l:�1hc��@m�#JN/� x��K�¿���#M��~�uM?[o��By��+.�j�C� � ��AEbG�Z�U�4�����^Pf��׮���6��q��A�V7V�:1��^��
�Qfmi��n��X���E%z���aj�|g��@D�(W�$kҶy-F��/I��5�6�Ϭ�0͓��C������ڻ�,�� �zu�m:�#h��f�v�]�A4l֋���tZT�6f�h�"
%+�LF�g�əA#k��-ՠDR�����&o ��W�K.�(U����jTv�\���;���'��vQ+�[e<����WCa�V+�|������C��%��B>O�a�R���$���g�=�b:Ӕ��}eRz젲q�Hg�tB�W�5�b;�q�F�w�\���]8owQBv:��0.�C���s`�[a*vI��-X����a�71oNՉ�B6E{Bn��t��1�8�*z�t���vL�Hf]��)�YmzU��m-gˠ�}=2�Ly�C�׬��n�X�N��������K�P�^���c`�.a�h c*��m�Y����k.��ٺG���׏�j��vy�e�MP9ә�fݞ�F2��&�t>������Y��B,cDו�nw[CԖ�R�L��#*ZY���sd�'��+y����(�%�,	�<�MH��л�W����f�A0UE��@(AU�/J�ʁ�tK��s�ސ�mOs�T�yR�����zn�60�~B���l�h���r���z
s�L��f,u��;k��kd�3��Բ8v^��9;6��8�uDɵ��6�D�}c��X��-��O����Q]���s�������j<,J�z�=�5�N%=i�?6B��U?���Î> ޻=�ɱ�~�R�"����(b��V��a�{|r.��K�ϋ��ч�M4��2Z&q:(��	��9࡚���5P
������n0.�w7�(Wt`ϫ