//-----------------------------------------------------------------------------
// UC Berkeley CS150
// Lab 0, Spring 2013
// Module: FA.v
// Desc: 1-bit Full Adder
//       You may only use structural verilog in this module.       
//-----------------------------------------------------------------------------
module FA(
    input A, B, Cin,
    output Sum, Cout
);
   // Structural verilog only!
   /********YOUR CODE HERE********/
   
   /********END CODE********/
endmodule

