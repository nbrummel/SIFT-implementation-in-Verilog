XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����i<ܥ�������|�>Ӭ��/�82#>��ď�
�������A8����.*�?��׆@�B"���[�,(���FɊiD�+q��7�#'�p�e�}����I�H������+?��u>zg����$��}S��ft&�M{۲.�V���]}��)Gy�p�S!QPA?����`
n%��1{K	�J��L���v�Dg�Nݻ�ו�9g���N��x����۟�sv�"s���$\o��+��M����h���ո~�;�����-l MG���,�Op�g�m�+uZ5�ɘ���l�
�we�T�b�'K�>^�	���7��L�����Z�u�QO����O����M�"Q�AųKØH�]X����l�~T
V��	�
���Χ�Ru���&�{<$>�_rcL��:1�ƧFy���G�.����^ư�DI��&�]B;������q#�r6���D0We$����3\�|�=z�2�".#����&��;���S+���L��R|�G��fՌ벦�#o�C_��W7������PҎ߼� ��	4��i��D��w|D,��`�[�Dx��	B6?���I�	�{���k�f��D�d�̛�+t޹!����ݕ�  z��28@��_p�8}1m��_�*;������
�K����p�g1��+��@Q�a g��E�w�%�y� z|{6x9C�9�,9����3|=��;�ݯ 4r&�>LJ�|m�r<s�,p0��Έ��s�6-��XlxVHYEB    2a4d     c10�>C��o���4V']�Ч̧H�"	2xV9�9A�ոG�w��A��鿉q�8/��pW�$s�V�4ά�|4�F�G!?��"#xa�bQq���i����R�\H�`��l\���6:�c܈�wr���_�]�.�oE辜����|ɻ�^Y��q���R`�g��b���^_�#O ؕCV�^��L)�ӿ؟\���7��-�Gb�!����j!�/���Y�>�`��s¾���B��,�=�r��x�/acyQZtKbj�k.��[��3˺�9kᚚ���	M�8�y��f����mc���F�5<�� >��H�e_�1I�.�]Z$8�֫b!���Gy I���uN����>(!�@��n$P����<U��b7փX������à	�]V�4'�`�FX2}�M�M!�xÒ�	O�v��#��s>�ү���l�&���'h�S�@�����v�o�ӓ�3�� �Ú|���7/�\Xw!����(�^��c��d�ڗ��z�ٲ�aP��:������s@��X��+�J��b6uz
��ّ׽��%��~�sp�!����c�����mo�� ���s�(�?'ʷe#�R%]p|����B������(��G�o��s4(�� Q� ���p]H�ټ3���PY>I�Jٶ�p�lx�9h?�n�PK���`���j6��Jv��["���aʗ=��H�����.2'>?l4_xx\�1��	��%E�(x���L�P��b� >"#��N3���m� ��l*��MB�+T}R@.Dz[$Y�?HK���z<핊&b�w8�>�O����g��V;D�6~�w���V�u?bcE�s�<�Hs.��6[]�7�!��.����ح���18&M��`�Bk�H�90�X�:���K��"�{)��9���~d�f�[�{ �����`���!M��F�3�k�	�ɾ,�:����#_Ƨ�\����jU˃�)�'�Maѐ��eJ{�7b8�!t���PO�e�ξ���9��N��V�����B����J�(6��xG���Q���=��nN�9}!�1UJR����5�):����fl��H����S����|6�R��@,�T\�,�l(Tӣ=
�0�7���Pp���	j\(1�`M����<2oZn��|;.�� ~&=�`ic�����4 �[g{�E�@����S5�z�����i�AVgdNq��،��yhH��P���9��뵫�iC��t���,}%O�8��|;HO������xMmS�Z?���id�gG��n�2��O�x�_;��t+��h�ޏ���^�\�j#>g�=�����@a����/�X1_���/E6N�+)1�ْK�W��OJ�w�v�ǧ�J�1*A�~:����h����3���l�иT�YqG���@��-��|k��of�E�����_9l 27�:���A+�#�U���t��
�X=lh�f�`�w�g��n�J�ߔ)Բ9��|�-]�xG��k��e���5�j;�1cK"��^W��Z.�#Ma��'23E���^�6_����*(����$��`�O��vk�w?�!�a�v�ĉ��-)�y��%_��TTq����oR��*nlο��%�	�0yv)����D����=�_D��Z��{��|��C��Ab,	��.�0���.^}���~�vd�Dƭ�2Q�e-(Q��k����i�ͣ�2��W%�5l��U��-��+\���*+���h+������OU+�g=���gQ��Q}�!�� Du���0��)�=�Ƒ|��.����%<��Tv�Eq��#��A��@��?�Y��c���{�j7���H��	yWأo{p�Ǌ�@U�I�˧�&l�&�_�nV��7S���
h����w�
$�u�(v���?!F�?�K�Ò;�Y�jh�Z��B�a�0�m��J'!�Q������!�^�����P4����HኅTD�9J84�A�˷(('��2�j�V�v��:�d�mk"���}"E��ӸD��&�0�t����1tZz�����q{\i��`�o|�V�4��Z�t݉�վ4)��2Z??ͽ0�$*7����xҔ�����t���K\R���W~��`���vZm�{Urh?�P6�C� 6�}9�Y��|4��4�B�zʰ�QLt�MA�`�[�AN�T��,��E'���oа��C�i!gy&8����>M����W)k�Ս>��cc�E۟���g�H�V߷��B�zK>�g���c���S��Bb�~��f�\!�N!�1�x6��U[�ԛox�:���h��) L0#�?t�vȉ����v  ���U���Q�h�{�ST��:�
���`ֈ��j�/ۄ�ボ�r5)v�*3�k[/���R�r��i �^~�ȱN�@�(��-2�g��]�E��dj��f�T�y�W�)�����',����?\��ln)�:��2J���~��tiX�4C�r�+=E�a��.�1��?^R}��Т1Ѳ�P�4���}��3�W���wY�{�T��w�j$���ZI`[�Nȍk#f�(ޠzx�T��PvͦeH��F��:�R0X��Q5H���鳏�X��Y�F��L���DY����"���5 3�ȁ�eGwz�ɏ��*g��$Y�8���&��x�A���/��09�?>^2���#5��S��Z�59S/l3��Ţb�L4�A��S�Fc��2`y�P�6����ܝEᖪ�����3p�,1'P왉S;�����t5��އ���|������R�Xc�>)�<��X��` ��ЅZ�Ă20"Px^�>�O�g�K#J�j���A(d�>D��λ?����oKhN�߄�7� ����V�_sbX���,Lѓ�H��ȖEf��Z̂-!��LH�$�Fg,5/#��(V!��0��Z%叓6� `�c\u_�Tp�$gT���
��=T��60�Vޞ�i�O�S
��#s�2^�Dp xd1��N+��Pu���
3 ������k`