XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Tq�E����9cXė~�> #�p���;$���.�5-����h(�^�S�S�?��R�����sT^�����$�%':�0E�IF�����H�h���	BSaD��s���g]w:z@'��J���m-<�ٜ]W��0c��J���"��< �������6��6T~��w�[��BI�a�C^3�M��5Y�[�5m��#B�*��9�F@Y�k8���I�����N�П�he]��ݒ�+M�����v�(�w���N?.ɾ*�����֨��G.D�qִ�a_����ӛ��.�pz�	���s����E���C]��17�/O�����P��N�PnP��&�-�6̻o�x�
<��ߓ�]�@Q/]8�ƏA�ui��*-R1��|�=w̼�~�)E�Aa���5e4�Nz�j~|Wy��tƧ����ʛ�u�����bB�B�[�~�8�Q��|`V�c��˭�k%ˤ�c)�3uN��($}�ݟ�P[%�I'�j��D�'\� �q��5�t�A�xq&o<-��Ar��z[~}�s���,i����V�E��JOf�i��9L��3�:� �7�3�:�)e?����G���a���y�$EL�r���g� �G`�����P.~�����q���ZF&PR���(6߱l�ů��h��"�i��Z�%��`�a�aP��Y���!��S4b<2Z��x���Y�nB�3�ٔ���m�R�2ˌy�:ӎ��0T,��]����1W -����h	�
XlxVHYEB    b631    1a00@H�q���*�׎9ЍSn����\��H��5v���m���Yc�d���D�T�6����4ϛ��K��T�?!�Ib[k�gէC��u˦x��p��	�}莏%}.ڧ���ck�B/����Mk�L������~�[���>e��48�+��+��q�y�{ga�o#a��������b�`z!7	�w�[� ���-*:g�P�����Y8�E>�t���\ �z&)]�m)r���]U,���t��:d�9L�D���YR��VT���4�K_h!ТUV�D�P�̑��l�ʤZ:�ע6�R-����[е�[	@�4$��s/�Z1=�;���o
�&�,�����2�Q��Āvu<JX��D*J�OX�6���|`���pZ����뒖̗�s$���߾y��қ��>�1�u���_��5o�G?Q��z��L ��ɠ5pm Ax� ��V�(�6�~�p`;���řF��YA��NzC�efGP�뎐5>����m{˧lbb��x@lݠ����v�0�AJq9��������*��mctG��҉:!���o��A�?�`c�pa��X&�W������C�y�Ȯ9I�Y�Q�Β��G�#��Fⴝt�}�������<-kC��wJ����6��t���N(�3?�i;i�
:��@���3-���5�U�E(���}~]�|P��L�ic��Jq�0ů��!�Y,{u��YZ�n��{�XR�)�05O�N�w��}(�o"�R�'|����tJv��ޮ$*�M��W[}�h(���S�e~�C�4��0wc�����
���	�+�����!�?SS=��������pA�Ѐ�o�1��o��wve����a�M;T2kh�f����}�^Z~*�`��q6kmZ5T�;�cSf�:����	���L7�]>P<,F
�S�*�s��9
��;�Ԇ��!�2�$9��5�;�o��Y`u�oB.(�L��>#���j���-�ׁ���X`�s\(X�|�·�E�р�2�mL�#B41"����?�S$.����9�#=��C�-C�t��+��T�xn�dd��rՏ}b��fs�p�1u���H=�q))�®Q��`brߪ����V��߹c@��^�$�����y��Y�fMɟG{�Y�`��
ݧ㵗|�~������٫��Lh��O<���A�7�(h1�zv�˽ A'y,4�lX#H���Y1�IӋ�k�����
4Q�o�7X�?e6���筕�����U��!x,�$PKu�7Ʒ���<t�/擽�KU	���d���Q�<'�"����Ј�#)�O�4p[e���8۷����Cc;D�Q����<�gQr'B d�����+C�T��<�@7]��,}V8����ΰU��"�<v��=�ɵ�f龝[�]%+l���������=�1��iY�L����ߖ~'fI�H�ȵ=�T����eR#z��0H�9ж�r�<Q&�OHp�@��>Kϰ@��7�eIX0�����<.?7�̮��͆��a�y��� $�o]x�ãTq�M�֥I����@��A� �m+W-8�B�AY�� �IU��D,��Y+b�lO�Ⱉۜ��
��o��m���b:�($5l�E�A�'����g�J6&3�ɰU����v��� ����V��g�t���%z.�5ֽ���0�5�����`�����[��=J�<��W�Ud�I�î������>x޾:(��G�/m���C�M�,Z�4�Z(��̎gg��02ל��LJa�mPE��/Y�u#���Nj��Oe��y��e��0K���!��Z�p��<=c�g�*'��ʫ�W��+��&��y� Ҙ�3�J���8�S�*}lP��~�0��s�z�T��SY<\�����P)\�����%G��5��v(�ǐ�y3n��O�A�JZ�T�&��5���/d@4�ƀ�����E�Q0ŵ	iu���4����`�4��$/��H�=���@*G6e�z�Iy���A�s����ڪp`1#��q#
��/�V��4��A��H`���e�0�M���@w1΍#������JH�-��f`G@x�VU�׎�����9�|=����\{儯]�C�x��F�lg�����Ĳ�V|���0�2�P����a �o�I�D�3;|��f��	!u���O(o�=��v�f~~ڣ��9�Ԍ�W�U����r"؉��Z���;��8? :���� f���K�� R��=όts�;|�:\j$!�����{����T�t��
:#y�L$)佋�Y�\�쿴xd���Ф��q��G�:	���:ӨƁ�O?�>���D�AU�m����=C;�p�$`����oO�<$�u�su��o2 �Kr�;Ώ���o�Vxht�`��[|y@*�Y>]Q�%a!��nG��<���F� �����J�DC�7
5�~Q�%'��c�vrVS}y�i��_d�0d���x�Q���=�%�$^HA}2��[VS��G�b��BTC�
����#�߯T�G�4�q*@O��ϲC+L��ğ��#�K �f{��~���&#���N�f;j}�)>����襨)��p@35	?$.z�oZ��L���(rvUXY
\����{v��W�4j
�=�ΝuqX�'N��H�o���'��� A�B�{[x��r/����G�:f1�BU�x���UZa�}GS�A ��X�~]˙�×Xd �O�Cz�IR�6�^2��0��a3G^~J����6�6 ݗF攘֣��^E�O|��os!U�!��_*:{���a@��(�ɧ�Lp.�}�ms�Ⱃ�d�ENt��Eȍ��w�AāA�Vb��%��&6<R�b$���O�y�L3U��"�ej/VE���yG�[qL���Js�|���:=`ڇ�ۂ
�d�W�k4�F��d���B�%\+�/6`r���˳���hS#�~�W;���>�%O���P�����L�8��^;X� S��<ɿS5����,���м����t�ϗ�AV�}�:�����s��@%�	���2YfBN�g�W�	�q|2iwS� �bË�p�Q��	�uq�k��,$�I������Y���E�s�Ͽ�_M�7����7���*5[���4����}]�`,�Z2^J"qZe_��<������eD��z����ah�Ϫ���u�^�|� ��?]�a9C�Oe|�A��.�dor1έ�[��^=�>0�`�Q�eL�4���(a����)��(c��V4u�c�Y�y���p���,��X"��4�(�)��)���U�T&{��%��w�K����$6���OG{�Ō~՟fd:�O�G�~.%X#���43֋����z)1�Kk �D��!�û��u�ˌ%_Dh�T���%��C�z��\ l����O� �c�v[��@,��g1��$�Ɨ�x<�0�2�69)j��ύ4�:�h{���0Mл���dHa6�<N/"�P�3<x�Y�C_W����������p53(Z��42���|M�=�ϔ�(�;Nwv&�L0/i���?�Y��:Ɉ�>F -�S���7��6�^�S,y����y&�Ŝr�'8��Ĕk P��{sP�W}U��r�*���ڣ�k��fXW��T�u��@���O� 듓���M�S+�,(Li�j-��&��Aw��na�	�ס0Kiĳ��-D4t!��C�P�Lӓ�fA�q�]L?�qZ�]��2�H�;SO)�Q�������ZW��PS�[�K�GW�V �+ZN����ֿ*��{�j�	]��d�>R�i3ƝzYӳ�x��J��V������-����Ҷ��3�;_��Ƃeo��KA�צ��KIw����jCL$��Ud!��ULqCL�:���&�Kn��%S`Eu��@�,g�QD]L �e8�mv<=^09�'C�Ǐ4�>����|�C�Q�2Ƹ��ѣ��}ԝ���?Z����
vs*_������y	ǵ,TcQ�u}��^�ۜ��T�K���>�/��˩�V7�i
���~��x�.b����;�����.������ �h�������Wz�+1���> 4��W���
�]��eR��<�ݹ+ܹmϪ�)$��O7����秪���:Ͻ���+#��+�t3׳їH������X��m�%(�o�,�`:Ȍ�3�s��_�]PIu������F�{'�� ;���״R��īw��;B�DŻI2`(�^�u؁��p��w�F�,$�/�j��3�g�bBHL����c{O�t���@T�B��#�r��hh������ �QE?t�'3g44�	��o��6).0kz�xR�Z��F0��	@2N�!)��nR��`��X�,N��H����5���by���0y��Z�v ���)�G�I�i����/a���ɡM@x@�a�W˅E�=���ŵ��t�-W�8���B�����y�˭$��)ɜ��L+z�E��Ñ�{j��	�YL�������6�R�
�d�o
�����j��s��r^����˓%��,Z
��������wK�Y뫮�N��T{��+��>J-��Z�" Uc��5識ĥ0�O�|�?W�l��8*��o�0G��9a��8�����xM7څڐ�C��	7E�0�?�m���:��0 se�W%j"Ob��3}g�{��"נ�Т4�6'��ÿ�'�J+��-ܴ �-�W���5i�p�WYN�����|J0��r&��=��vLG��Y�-�p:C	
"�a �dl�FE�8�%�����5�f*B�<�<���.���9����Z���CO�?%
��u�e>6�Q�4�����]g��W�_��M����]����)���<�څɋ[�48�Em�Z����}�\�+�.��1v>R`�N��+�Ab���34�����"R�z��v�dZ�,����t��$~Ϯ����k/���]�6T�\�`��*�i|���?�����E�kӈ��S��<��D��_��~n�8�$5��v0�%z�ۖ2�������+. �E/9��1	�el�n��9M��j��y��Zq����妁��l UG[ �l�,¯�QW�91�4RN��ֳ�([8�!"�����I@{* ���2X$^�{�e6��y�Q�eC��K4lA�5��܁����-v;�C\|���BL ��e�����������˩�HK�&٨5�bX#�y}̭�C�C�/DE�����(�w����7UH��uvx�sw<Ζp+���t%�θ2S�j���A&�ع0�ץ��84$�u�	�7"�:����_�NѾ1m,tfb����)����_c��Mvgp��W�l.e�<��e(��e�-i+1��۟`�ʯ\��3�$����&���^`����I�BT���ɍ�)2/��k\�����Oe�ƥ��1���mh�;�$Kp^��xJ�JCy��^�Z17�Nn>F:o���4؃h���u�jl�.���$5�}П~�PI���SyEG�v�5�rϚ?|~�CUD��ľG��Mn�����uFz[�����˜n��m�����MT(|Z^�� >Ն��p�|m	/ F_���`��mŜ}�-i3B�ڗ��e�H"h��-�ؠ,.������:��p��?���=75y�dY%g�M�i�y�z)�$]p�S�LǟI3��۰I��g�I�WOs��G���*�z����m�ZM���P�<W	��}ݬ6��{dw'R��X�zJDR~�6_���S,�	&R?z��AbF�{������ެ�{p��6�ѫ8��A.޼ (M���Rp(w��!D0N�����c�$D]p�;�T��袿!��G�q�C���DLd �Z����ȁ�&���&g-�n����eu.��\rś�G�0_eyP�a*>���'F��7B��������2����2�&-�i3�-�ҩ�K��F�X�������n�ӷ�kW�0��aX��	���ZjW���;Oë�E�zCTo�-v��/:j�x�р����\@��1]A?�;�^`�rw`H�Y޳99!*���3uv]�V^%�Ӕ�&N���}�?�G��e|�W�e�9im���������G�km�	�x���/�M$�ꮙ�F�����ՋB��vT�:��b�1��w��Q������E0���C�X�0%i��.�����n�|n��d�k�}a%#M� ��)�5���ݬh��;c�Q�y;�&�+S69�q١�e�g�:Q� �6D?L�k�lxEP\���@'"��~���a|�s[s��Z+��Y4ݥˀ�=5�}��?�;Z�����]C"Iȯa�V��2ޱS�_A�]�YG��?z�qܜ<P���-r7v3}����n�p:?���oMR:�j���!������C��n���Ǒ�m���*�}+c=;�N�C��Ƽ��_cAN2e���� �#Q&��YOQ�c�i���1PrB)��e��Rc� T.��s�->g��^�90\�]�pAɎԧ��>��҄�!?�i�틄9�\m�!H��ՖO��6�6lew�%Cm*'�