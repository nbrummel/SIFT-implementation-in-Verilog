XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y�1�rw�[���Z+�E�5�D8l
�{\�z���{kM��A�1	��h�Q���4��Z���nH��X=ص� ��Mt-����MJ�3D��_;���P��y�`��Y��P!`�:sz�K�QG�[�kܡ���N�Ԝ)��z��d=�E�=�jw�ߣ�7)˕�*�ٖV�s��eX�5���k3�\8����C�����M���ߥE�Ü-��a+�.z�v@��h�<4���
�����֧����^�1��[hI=���ǚ�����]�3Cz�,`�C���n����n��q�.��6��u9\��	{��$-p��\̧!���1�����g��E�9O�I�I�]���N�N��Nq=�����*A�����H{��G�_PqN�Gz�J�S�;���T�a&8�H=��y�?���w��X�X� ��i����`�7�@��[?�����#�ȵ�=LLY�����a�REe��K���UO�#�n��,�s�/
��U��[F���GCzTG�e"4��M�Oz�V!�����	��;��:���P�q��!)@$'h՟zt���XhBk�h�&M��g� �E���b�=�q0f3p�fgq_8'���+m�4�y��������i��٠�W$�M{����?G�i�'��52� ��(OX�����:��I�\u���g�_v�Z�%��I՟6�� ��OCKX[D��='��]2=kU�6W�i�H�]>�v�������6�:D%�j�XlxVHYEB    47e6    10b0��4�[E/"����a�Nu_�GxU���J@؉b �Sv��X,�$J�F��b̑����o��Ɩ�yg~b���D4z�mC`�v�!�с��Yټ�
"z�!�ך�+�x����	tB��|�J����#�
�}����H��hW���Ke�����/8$��|R���\�\Th�3�=��?=�4���ݾ5������")���$mJl����-[����c�}+&?�Phw?�Z�K��`tf�3�6�#ھ�WP7��ha;4s�?b��QU�������d�u�;F��V�iǉ��/�}�]�x\�'�1`X@/sUk�ǲHd�ĺ1."�{3Z�;���1B�9ē�#\J���m��u�"��z#�W�7��ܡ.�ӑ,�����uG��%�����j�m+�����5�q[+sΝ	�U��+AU�(\.;@��N7�0�<��ۢ�c��4�=3�z�Η,t�ʛ��������B\5�����򕚫7&�^��p�N�Q3H���#3��a"����dN���@���m�j$M	d����B�ﱁ�*̵�n���<�4������~N�@Vg2����E��s|�' ���ڨ�lG���ٟ~���V��Z���t�N�a�%|i(@z���b/dC��Y���7����I��"��N��h�
�l�HR�K@�\��Wb�X�m�9��kȤ@��+ߞ�hU�	?���;�7��9/m�������������b A1%|�hmH�Atd�{�2?�!@sU�Ctq�9�R~���\4���� ���?t�Y	�!
z)E��6~���^�&��~E2�������˒�xr�y����s��t��Z��]��"%>��i��c�V|�I���Gq�7[���	�a�%E����j�N]��X�U~f�q��,`�|��"qm����f-��3r�nlM�uz�7���:3�?�nv��z�p�P�+"��������!v08�Z�1�!0��=|��S�������f���o�'o R&EI�tz���JѝO�&)�ǱM�O�vW�¶���X���jBn��5b��E#p�O%Jk�x}$��d������ӟ���U����ϣ�!��F�b�5f�@��r�W�H_�D��&&$Y�!�04�d(�YQ.ۃ�8($�P(�9��i"�)U��;!!�7��)_S<�)SA� ��$�Ӂ5���k�aTC㛵p�K���(0�CY�|Rd[d�ϤZ,v����ga@�`R���?�:Q�<�*�5��ư����e������S-���ND/J��!�S�E�h�`���X嚁!�,h�k.��_j�}v/�?.Ls�B�КZ��ƈ�]N�����T����Ns�ȧ�8`���(�Q�F����>u?,�Y���33fiieR6oOct&����}�� JE���n}0�?E3��`e���:���8���/���w�r���w� ������w�;x4��H��.���TW����!(ZL��i6b��
�o�� Ha�>N�mNXU�pQRa��P	D,�Ͼ{(Q�O��e���Kn��H�D���xmMM�U�c����
Y���%��%�~�Έ�v��b�Bj�V��d�B�x(P��"ىHW�,1�쭣�ɉV*��Ug:� ��v���'��e����B'�+���F}RöK\}�E��9Ԃ��:�7�`>��G��xU�r�S]��t�����lwR��+���eO�?��A��]� CG���&��r��Z����'�	��3(kŠ/ZV�6�A�	�x�[,�p_��Y�5t��=(����0��7Q�vҘ`(x4R9[0^����c�#R�!�\-�Z|����k��/�Jj��.�!cN怑�G
;'�HW,8P؛¡T��H�f��5�� d����O���w��[�!X�Y���H��ILÉ�&�lG��g�� %��錊��/�0��أ��z����\��x�~�"����M{�:R�9#�8]oy\��@�6 *�M����{3GQ	��lx�a�d��u^j��
_��17�{us��E��~�K�)dt w�AR���
���׵{�����1N��HW��p�Ϭ<�wc�d��te3_�$�{�?#����y�*�6�Oo�]0w�8Ә�#�A|U�]%U�����j�pKHg1m�$��Ž/9��}�Z��ު� ?S�Eڞ�Fk��:�̣Og��/�~?2�৞�]�oծ!��u�F$:ր�v@�e��Q����&a�/E5]k��@���8+�Z�54�8Tk_U���r�sv�*�D�f'�ǔ�$���A�HA�R�Ds��
19+�E�.O���7���_u?C��	g��"�H/U}�2����G�;�]�|��v�u&V��	a�US��p������d�)㴧��$�o�\a����;R�3����-`f�{�/���p�lU`|q�'�.� ��[����_�@������GUlO�jV�b�.^c��БT�J�f����{�J�[|&����Qd K� a�X���B�h��A��j��A���ǵ��=L�L�8��$o��	(���a����q���H}l/�&}j��n��~�d�a�lJl�~���ऋ[�/	�u�������J���}_�A*�DO(C��%�8��@@l���<2_	��j܂(�֗",T���+��Գw1	5?}u�R�bΎ�5A��B��8���I���Hqpˀ7��uj�&����_K�y�N#�	�+J��5����b�t�v�Y����_佻��֙|�m�w}F��������ٖ��򛑫GԊ焆��	Ү(���8��Q<S���jr�z]&ҁ�w��+i:y����� 0���z��)��Ϣ<�E Fc��״�Č	ĺ��RyY��r��b�9!��&�%qw��U�9�����Vh<92 �wV���ܲպ��`�����_�opz���h8�
L��e����x�,�,[�Ucp�O����ǎv��Y�B��~�L�/e�iS��]�伫�_Nzry���l��c��4@Q"���⭀��"w�_F���6QAD)s����p���DPz�e �"��,9&*?�����[���# P��[-AoК��4��L��	&��1A�����~���s������ٽ�V�b��v��_a�'��#m�k������ ����J)Ve��Bq�m�q��a�cܑ�qi���:���Ϳ��#�,s����BAX�hV�e+J����t][��^����C��Gǌ�rԛ����u�B��l���:�+�)�x��\�^l&v������5ʆ"��l�6f"�5��$Uy���,�d�E^�F{W|^~
���Zҋ�<����Nt��7<�t�zoI>�2uR�vk����<5�������7�:����i���3FQ�^_�i�0�k�.�����Ġ����Pqb���.BX���7*�u,����Uo�����<���1�X����tZ��b��I?�s����.`��םg���+^ 8+]�&
�����v�Vt�Y��'�D�*�Q���1��C~����}H~ʺ;%X�.c�;�kAmT�>����f\�h\���Ў�@�̖�C��:�8���N���[ ��Ty���0Ֆzߴ2@��L/L�l���D:4�'�X&�����V�5Q�WSP�A�.��Ұ���'ϕ�2ᵲ$�7� ``�#ɝ��}^vP�\L\3(�0VT�	g��^HEVz��
v]�=�~�9�v=�k(�r�	�{(�)���|�\�`�!����K����6B��;��1�}fĽa���&:i8!���z���:�,��!��%������D0��E_֋��G��=pe�:T-�� ��A�|x�C8��UW�t%i՛�	1�Z/��l���^�>�«	����O��m��@u,<�Ղ�H�ax�gA�?CUK\@6z������Ht�%��'��k���2�JsZH�Sig�2y5=�CY�u�_F���q-���Fm A�����t�����S͸դ���;��y99M�Ҟ<�L��.������;\2��"Ҩ����:���� ~�3��z0���12C�>i��C�!��^��U�D�@n�����*�ȱ=R�Y[ě8�W��BJg��v8���fL��e��ϡ`��曌�	��0"�6���C�MO.�k&����U