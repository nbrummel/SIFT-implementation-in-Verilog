XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`H]}�7>' ��=t-�)>\�,h��maI�W8=xLհ��{� �,�_?��|"�3����P��QD�
��%�ڿ�����f"���B4�����P�!�`go���p3�G�i��B����@��k�n�-��讘1����-R���Mcp"[�mJ�D��J~�ױ	�a���)X"V`A�K�`�c/34�_�֥-l/<�l&�P�g\\�����*7\'+��hnX��(c��y>�����D,����ŗ	8 ��.$�����0ԖDJf#8$��/N#W7�?��]?�eXmT�3"=p�0M	��'�eZ�����Qd`��ڴT�-��
p��=AM�?�L'��lS>O��+�亟�L��U?g���	����d��L\�;f�(�."s���b���T[÷Υ/�L9��y���a��p���a��AL,�<'Gl�3�#b��SR͙�*��ɇm�2�1jK_��~����O�VL�g�8�wW�M���V
lg���,ǅ�_�cq/��3��&�,�t� �e�d��W;d���uq>�P��2��oXKVRY-8�l���m8��RF�h����r��y���%�7��s=�P�+�!����<���}hx�·�ò	�]\�6E�	C���!�����2�oI�s�r�X2�a�TӇ2*�6�%�i�E���0��Ѹ��a�yI���UA���&(~�H\wS��	������T ����`Z`Կ8�ڱ�ж",��~�X�Y�N�5����D�XlxVHYEB    6610    12d0�0Sޓ�� ao��H'�7�e��A�8�&f�'4��=lɡ	�mf��(�Zc��4$]|UJ���Z�k�Y�V�
M��3/�(��[x�Z�*������|���Ј"¤�M姿}���)��� vp�|�+?Dm��ȚO�j�h�Ti~UH���d<F��sM}pԸd�{���MO�L�,~x�@?i��3ah�� ��i��U���iNs\}F���d��%C�����>�M3��ߙјO�lnh߬��c�G�����>��H��u�|�W�X�1Yn��\���2��A,�\�O���y��6�r��h��2iL@�0s��2d7��!"�3�];�>��)(���k6���D����0���e܉�6ϋ�C�Gj�Uz��C�,�ش����q=z0��|�JǓ(��9(�'�e�@�C2pFh�y�c?�R�e�;1x�|�k\{��J��~��D�4��� ��BP�;;�e(|�q��;�'�J��aN|�R�L��J�0;�Ʀʗ'jp�����;��v���¤Mwڙ���6�C�U��lbѳ�p6y��ܮ8�-,��k��r&����W$�_�T����:������7}�l�<��W���{�D���B�ӡ�M�Cm<��W6������6�D�sԯ�yH�b��Oc/��P���b���5tgwr�;���;Z�3Y>���w��Nh�s�Bhw��L���"��9�PD����0�P����G�޵A�lJ����h���g�s_�� �Ģ�AD⬙Ňz������;�Ƹ����5���j1��֒!*
�O	s����mΣ�YeI�v\�<~�=̇�*&7C�^Ύ�g[?���z Sa�[�����A4�������k���v��+-˫���\U�� �]�[��>e���d�	ۼ�*զ>����P;��"J�� �
g��o!Y�4�71T�Z����Y,�ǚ�1�GxDg�o�nV��rvuL�o���X��?>H�iSAL+&�x^r�H��g�){�w�)A�.:�9եs+����\m�&߯%��� �c^l#���ӴN���.�m�:5�+q�:*vf�b��x�o9`ɀ��'��^�j���?�_���0�ۉ G⥘Vۜ��%��iR�b�o�2�II�M����t�9�d6|����⸰XLJ�)z��&��],�~�u�(�l��ۑ��_(�����G�������gO\c�ה�0dv�P��H�[��(����?�gxq��d`x�O�����4*@@�]NUŽ��d��~r�� U!Q,�+�	��'�zYAqr����D<�C��i�D�d��H�4���}�,�������ǜ����?� ч�f�FS���l���J�hSx�U]Z���E���HN�c�&Y�kY��S�fiz>�yB���
i�.���!ꬺ�y������-PP�Y���N~�6����l8L��w��;����vL�ElW������j�qcNڔm�ӗ��X:����ׅ8w�P�������E�"�'�De����%��诸���φL��_~D�?\�-���R_(�cFvn�i�����4�
^}�"T�	,C�	h��p��� �J|�ì�/��{�מ�Ɠj��
y�C�q�R���4��723�!�u*$~�T�&z�������r>�2�]�����.��V(�U������o�Dᖔ��{k�;Œ���v 2v� �@�WU�cb0Ҡx�`r,l���c&seU�FZ�oȑ��$Ԙ�n�/��!(x`Y@�q	��($I2�,�|
��A6Eƨ3�7��M�fH��9yD ��fIU�N��0B(:o0w&�ۧG�"Λ�v�2s�La�=T	!�P�\��)�*/#��R��,��p~.;L����c�+:��?g�5�UF��؃&@z����-[�'1��̊ ��q�ɴ�2qbE��#l�Op���r>Pc>*���;V���K�{��$�d�Z�>���fZu��J)R��"�U��Ŭ�# �hH=�8�#p�gK�/���wSOk,��딲d�hn0[�+[\{ɜ�~<��B~TI��{ ��_Zj���h@,�q�L�6Bo�ɼ����1�+�y�+�t���6�D��\)�D��
��	��2T��(���={ˆ刑�U�ş��:�7���,�O�ϥ]�mM�:D���*�[O٣:��(�+rh뜲k� �H�tZ�����TCZA��:�Ў<��4�0���oL���zy�Pt=��ݦ, ����G������ի��.����`�Yָ��%r�bx:�*\h1�I�M�I��@:Z��C,Hx��b��1�0�إ��@0C�)��/�n_lTꜾ�|ԙ�Ì#��X���Ѵk���=���[�J������h{%����Fn��pZkǜ][�gBU:VQ���7���4f�j&����-���Ѕi ����ⶓ�r���N�[�sp�)�iX��h�x��a��ٹ6A5�M��4�H�8�r%�x7�h%�� �������a@�}߱$�;�9��@ʲ��:�b�SKo汍�����Ϟ��m�b@���uՑ��#g��?�ֹersG~<71Yݒ��[شv@<i�3��gF��,�}��#N�gـ�w
D�5������2�}�#V~2�-Fe	%v����Z�ʣ�O	h�^�"�%��cr�4#��v���8�}؇�5뱢�<S�6�O~��zM�#�v<S!�h�=r��p�_7jS��	�W�O�P#`n�(`��k&r��}��M�U�/ST�-�z���
�/r�}�cԹ	�qt�r������e��n���ɨeKc��"��]��`EH��k�h�ن�5Ϸ���G������l�ߒ�O��w���������;5RDx��W=���=�p��"�s*j�����d*|$Py	�Ҷ�,xq]�
iFMZ.�ρ�����-|�5>>me��'�<��:i�K^� �~�j
��N�7�+.��nK&�ց�}�� ���s�:�N-�k�8n�ǁ, d���7-�r�)��� �����%���� w^F���|�Q���=7�B�G�b7[�8i	OH~k�[�;��������e�N�� �Դ�!����@[g.�a��%?8Cf��q��(�#�$���[��i�e��R�1�֥5�ё	���``IbX��%r�	�G�]Q=.W�H�+<v[�*b>�S[�\/jDJ�}*�� ����OPߪ�Y�-�ĬM ��f����b�=�x0z�>K1��>g�s2. �.n*���
��]X�����#n�I�����i��p%t�o�I�,�5�Sb��ö���q�h����M�^��2M��Ѹ�$��E�p15%E�>��{��?�r�Փ��8#��2MW�I3���u�����ט���Bŗ9�ʂ���Ɍ?�I��쑹DÝ��U��ʟ矸D�j��EIw���F'*�v@N�?8Z�g�#5�L!O��*�{օ|K{gI�4�&LʷXq���
�����5�����"^�5);uPp|ȗ��\��qs�,C�������8�B�����{��#G� -�;#)�/˦ǡ漈��9�}2�KH% �S��GE�gׄ��S�� ��OFb���S��k$���oU�˯�ڬ�;oRg�2h�b:�ڻW�!��o�,C#�<�`q(�?���n�V�>:�O�$v��T���}h�v�u[;�����O�L
]#@U5W�
�{�(��/6���=3H�Ң�f]5O�6����3њ6���3[o�cÂ�}��a�b���?�N�M�H�21u�����0$rkapS`�W�͛�	�Y�YD�|�'��%��='\;)���e/�f!���#`GY���R���?���#	#�1�_ei�R8�D�j��"��������͏�E�8>��
�&�}6�+ɞED�w���>��|�(� G~�Y��T����-Z�Gɯ��&��8A��al������p��XA��g��n�O�ۥ"��ֲ�1|�(-E���r�H8�B��TQD��ݫ�NX�E�їf�q|�f�a:���r��l�>���1�X��S{_Ŭ�7u62�<��I�96�ܱr9\�۹�K7��V���|4��?�i�Ԇ�t��i���!���@3�'hY�>�'n��Žغ��!�Zc��҉����H{�G>���7iM�%��l�E(�zW��|�kaX�2-�^���#6z
���sf�k�`��${Pζ�&p����'99��^��Cݧ��Ś��%�-��t~$K��J��ң���l
�WOS�r�?��������V"%�X�<Ivr�����ۧ�S��'� �1�F� ��1������P�	��m��އk�2ܿ,��K� "q��6�2傞�T�*r?�ƄY%,�*�h�R!�z��{��0*�w4�@ÓdJ��A2���d����* �r�	��u�QS�R��p�lE���]�
���9�t@O�o~�g7ч7M��Z�Ĵ�	��������TV`:�Lz���m�u���v>�#���-ii��-ҝ� ,L�2�ە��_<�}�.��ﹳ���0�y���	e�B���s|���Y��څb�C�ʮʉ:�j�/伋�y?���LՌ��N��������W*��j	DI!����>���Nc�F����ќ|xg]JW��z����+1��懢�-"�x��.L9 z9C2��hԈ