XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����e��b��Nt1�� +���B�8cFR��S�6ꖾ{���}�J�i�&��$/�T2Y�G"��ׁ�L'���T�)j*���r ����xԀ�P��,(݀������R��i�{?��jD��)�����P�L�:I�v/�皕㔧�MlB���2���eT��"MXRF�^j_��&�F�{�^��nf+����7�B��L$��b,��ٳ:��!��[����:�rq��K�gٕ�����V\�2�h�� 8^�<ɥ�����U�v�R
�`uw�v\��x�	� �Lü�#c'Mzݵ��۴I�2�ţ��J%��^j����w��'�z�f�Z���U�ϓ�g���[6�@\������:p���kF�Hwy�f��G��'�7�0��z+M��LE���Vw��w��|W v�do��(h3�!�1�
L͠�`��,����Ǝ�wYmNq��Óu�)d��F����$G�f��:��Wc��P���ojK�B*p�BB���Ӈ�OU=9�p���n�o�jh�[���pX{� $�?i]�D�`T@��F�X��H�oH�]|j��D���XX�	���H��WV6*1:*�������2-Pb {��Ô��#�WA�	��2:S��۩�`��-_U�� Ѝ��-Q{Ӯ��6�(-���l�,C�����Ҧ�aW�;D���;�%�ٮ\���?:bq�ҕ	���Sřv٭Q�>L!q=��A�]�r����Y�<����p\ҍ��w��i��dAXlxVHYEB    fa00    1fd0�QPA(�xǭ�b�� �Z�{�D��7����ނ�}�/ ����4�( �3[N������Y��}��!?/��F�W����� A�R ,̝�Zp�=BS�+V�.4K�H�R���{�N����ø�8D������l���������m���uL��o����*3��|��U���)��fܖ��@^7c���!����:��+.Cd��lE��"t��r�A�_����5Bo����/6�* +���pSS|�%򶫿�O�)B������a�Y>*T?��[v
pT �Ͼ�ѡ���ÿD��	~��2�8	�fP���C�r�H���x��Ȉ�� ���i�9�5	���.����G���(�:�#̧��Ӎ�@	�U��Қ~b�V����>"���=7T�Q��]mԱ���<��hGuC�Q�Z�*������K,��q��
A|[7�gݠ ew���n�o���ZJ"ޜ�6w�uCR�t1t�����*75������ ����KS�=K�p�։���Ф�5����h#Y�;ǆ��e��<��j`�56��((�1�X[�����`�)�h�a�����<���N�T �ڣ���
v�VZ��8��z{|$S�"�nF��|Y�8��?�ET�U�)3�������&'ʎ��� ���0��F���7~����T �"�}�58�#e>(����\��ԛMS	����Tx��){������@�h:J"`��q�I�8���*SaH*�lP���ֽ��B�]S `Q��=��^�bg�?����w�j� �N�B1��Hj�P�d��td]c�;L[��5���u�]�|��x��ʧo=� `p҇{#�����.�t�!����(�ny�*�n����d�r����
��o8[4�~>S���x��i�	�[ޟ�Fv��?Kˀ�S"���{n��e�o'�2�{��Ydҍ)�P����؋���nm4�M,�4Y,`W%�>�� ��R�6y�H}��)p��qΎ�۪1<��L��0E��7l-p5�#�wE�XG�t��ѐ$C�6���m��Nm��+�x�T�i<\�?����CC���8�����ٞ��|/,��;��D,���P/�:��ܺ�#G|�vg)� �xs�� �_a2��B��}ޘ�������X�PBiÆo�5�D��l�*:st��קY�@���A)r#5�vh$�Y;,��m��,��̨�U�u� 	[�(���9z�,�s� %+VAb��\B��$?�JoBvr\+��~���P�w�r�G+.�Q�Hr�pF�޵P��^x�������ύ�Ǜ��2>�������{�z�s<hħ������txQyL��!��snL�*`����MBv4֧!PGب� �{�b=%:��ѳEI�1$��/YDq�_�B���cRU{u�lx���Gp���`���L�Y����<�Y��\,�T��R0�R��NŨ�}G�?WዕҎ�^�_G�UDS���_=��+zH�?#�mw��&Y�$�����J�DD9]U�4�>DB�(��4`E@�/ad����;@���螶�K�n�g�	E��5V��kT�g���o����V2S;�އ�x��u�F�+YQP�MlS@�W���7%�K�}�?Ս�k��7-���kK�=;��H���>d�<�72�����Q�>`m�w��c�U>��*L6�R���d������^�.>����B����2��2���bË��&J+�V"�㗽Q� d�����}/���
h���2ItC}ɒטCYbVJ?��I�4�X��fh!.*��j��-7Wȣ>�,�AC��\5
E��;~,�fW��=�H��ۨx���)΢]�&'�~�]T>^w�g�}bI��bI|�F�3�d�!>z����M��g����z��l>3���Y��{ �$���7ѻq�7�٬l�������!�oYT�2�.F�,RO��h�-���q[�L��-�QJɸDXW��U��M.��7#$�= ���&զ;}Gz��:u/�|�UObd��8�MfXsؾ���Ҽ���9Ά��U�M>Zȫ\��	F�[-�����	�p���4���1�J^{��k`z^�b�OYV?mϡ��Rײߗ��?:HWڂ���f�)�fk;��Mj���0�!E0q�{b΄}m�������q֑��a#�����Ƀ�UY`�P~\Q���t?75�r�����x^��yK�z�['��+F�M���>>u�J5�K����¨��Jb�<֋�
�@5��0e���r�DW�\��9�F��g�$�ؘ)��h�����Y��K��r��wk���g;�ݣ,8���J_�o0��Pi�Xͧg�R��c"�XK��d�����A4O���%X:F):f����^^ͽ���X8�g���I[}�z}?�9�1ñ�O��Z՝��(
|D�:�Jm��&>XP�,
�֑�oc;d�,H﨏���9�z��.S���O��,N'T���`-ou���>����=�̩��d��ⷵ�?�ӥ�d��zh�"؛��[��]
�|ڝ*S��w��2ņ�(��1��@{�a�Hl�|*�s�J=b�Ɖ#'��J0��w��������"�1����
4�I���U��W���(�� ��%��]��B��"X5�9�l�0�Њ�&L�e����p֟���#I�\3_݅F�ZOء�8�b�Ls��\jr݉�/,�caf��7(7e(�cz4U�eT�@��9��4���Q�<P�n��~`�Hߡ��2^,�Z�C�z���T��"[�.[��\��g:��}����	�L���5J�9��&w
B:rupdh�=��)��|]�8p��	�Sn|����7�=C�g�k��1���Oq+ m1���!���x^wKb�(0��U�`$��u�jnó<\}�oP���*e���߿t��9�x��r1nr�O���7'"��J�4Y��.t�i
�Ƚviņ��tā�O�a�}x�-�EּS�����������F2��^Ҝ9���$����WU\Աy��_*���i��<<�B�����y���Pv9��N��I�#Wp-l̬��2�=jбø�E��=�z����l�^�D�f�[�*�ǚ?����Z����>2�L�y�f�V��(���")V��T.��L
}p���r;���S�ڌep.#��1���u���(�C\�j0�R��\6�*
r��j��=k��w/��ai��b@�,�\�3q]r,b8���D��C?���:uʲV���j����� ��(���Px��n�7�G����KE��^n6SZ	`��"eLTj����a�=;������Y�"Vղ9����[y�Z?��5��3r�_"��ʍn鐨Y9ſ4��Nb�?���If޵��s.ж��� ��P��r�:f��v�
MA��̘B��"�)��#<�Ba#��{4���l� �h�f���+�X�5�v�yS�d�e��
��۳�v��j{����6�aǊ�����w�� y�5
ޞ�9�>�� �pyeiL)���M�.*5^s|쬨&��Xk�u�#����+�5'o�Z�<����dY�zG�z�{g��? ����o������[��7�a�%���u��ӿ�8�4ז�Oz��K�u���/q���w��G�&8 ֊�v;��T�Z�,���_a�%��-���̝�!�Ty�PAqX�gp��I�N�5
�R���S�J�}�8�%����ގ�w{�~MI�@�9�e�8��+H��y(��/A��WB�?�E�#a&:�}�8�n��F�Xʜ����Z��2��±O�rL��N��� m��#_��Ly{,C�%��\Y(��6��3D+�� ��1�nR���Q
�R����S�x�4 :�_ԇ���z��'|W}��)kcFe���v'4�ʇ|��d�rh+�^�?~��h�  ��13��<�d5��P�ɺR�i6�K������<��;��}����_����%�4��S<0���B������>s�]��4]4HXxT��6����V�S�Ǒ'X�R!E*N��æ%���6.��6�%Bw#���dz�D� �� �����7BK�7cl����$7v�,[�]���K��՚�������fVv ,�	B�ѱe��\].rz�5�f�ua�&,r���� d��@N������4�k�J��%�"�@�'��{,gxz�\�k��O�U2�T��1��ߟC�"��U�#��c��:��|�h*�!Y7Ջ� ({�%�y����
�l�n�/��`�8�q`���"��H��'�ޕvY���>}'ҫ��^*֏��&*�6���J�E$�pS�nA�jV��)���=�+�?�+�*P.�Y.�ѩ�F��z�{�f�@�W��Xh���9�zNn�ŋ(AZC�-������/�ȳ.�2j<R*G]�G�D[��u���Ñ�h���m뇷Դ�H|N�ʾ�Sw�:N���q��xg�w����RCvB�������9�i}��r�D.�Ձ�O�:xw���0�� #�4�^�0h��%�
�G4hJU�/�d�j,���(T�9��	�s�#$�cū�t����o˼<�5��^�]���������n��j���_*�@���xY7�������M�#Dx^�z��e�}�}K���[ᛱ�'��5�2S?K�eE�2�[�bM���<�2 ���cw)ה�)�|H���R9uKI��/� Ǵ`r���%&:�-����M����S1���z�bU��g��*f��"�d4��;����Y���D��O�E�M��/��]f�AF@��&��*O����J}��G����;_7_��x_�ma�|��w����,� ����VR�>���(c��%~�l�⎂cU���p]+ŋ�>�D���.`�f�����3Z��!h��C�W:�ک���@ڻ��4��� �X0fH��@Lv��|�h�V(�<Çbo?'�~���Pz���l����Ł���V�m_�Gx���t..��ׇ�Z/-LJ�{ם�Β��[�a\�	���l�������^}{3Q�x%G��dj�ֱ�1��n8�Q��/��s�|	e��t������J^I߃�Rq	Rg�S�[� O�(�~�=��G�偿��^>��f���I1�j ��G��V��fΊ5tIS�}ٶ�`��-���Wa��	�q2g�_rC�fGz�J����2ں��|a��M3wa尠�o��f��5�x�)�> �_
rZ'�8u���6�&���BrS���㹟f�wD�,�nkv�Df�{s�Xr)����<��NiW��\a$�{8\�$�35H��4�&�X�?����u1о=t*�����p�C�B�+y$;�	�xf�/8,=���m�M���I�������_�^	��u���G���g�Y�|0q�ZH^��m��3��d���Ǳ�# �B�"(�S��dA3�Օ��V.ޤ&����Q�2m�F��b	����Q��㮄-x�||=!��h`��
�%�5�M+c娨�b# %`���p0��CGyhdv�>�L1^�2}z���խ��|/�c�2���`8	����"���YCM��)�����ˮ�-�;3q� ��*#���Z]���5�!	��7�a$yٝ(ʷk�v�L)Z��gx�\�ě뷈i>�v'���y��>�H��&�v��^�s$�Z���QslB�3.*E�v�g�h���5Qzۢ���,Ց�@4����d�<�����4x���OWn13j^Eo��C|�k'}y�}԰~����୤o�9��L��4�EdԷպ�T�s4��W���ݟ�}|>�Z�X�D�zQ�s�Z�.�MO��>2q����_e	����-��dY���-������.Fh��Q)Xv)���f4N aU[R�N84H�ޙ��v�Y���Nt��j�$䮐Zp�ɂq�'�ե/��b��q��@�A�v�y������Dln�ULc�	U �3��{*Yr�?��2���$Z�LѦ|�YT�D�)���9��h뮄��e3L&�~�NW��p��#k�{�C-l����R@�h��NDln��󾑎xҸ�*��''��ы-�Z�{�[>�	C�c��}�tݛh�"��)����&oe�$Z����H;��1ŋ00 ������N�?!5��Mӳ��^����0�����z%r�m�I��Rmu�zě)=�Q-��p݈��
�V{3�a�盗k�E��B�Ë.K=f8~/�`%��k�V(&���Z������I�A��p�X��n�ζ���F��]���d��/*���!`>셻ې�cA�TWr�W�+a���1ɂ�ܤ���W��½Ъ���A�	�]]�ɜ��~�P�
��M��jÆ,��4�-�@��!����`�J��'K'�X���W��$g�x���NP���C�rĊ��i7ꈱ-��c�'���PM`�ܑ����ȇi��j���*-�%�8��Q%��o�p���aҍMX��� "�0{�����/�����ܡ�|+�Y��}YV�
��R�Cnn��o\���}F9��D��nRJ-Dw�6��6'K�c?�[ń�3S@~Xjա�r���SXh�%�p��~"�QW=l�p��$��X�;�C����o����f?x� j[�'N��(砧���
�F�Tȡ�s�C�c�8F�Iyz��m��UJ�O� �un��*lq5�-[�d{�� ��_���+��޾tP�4�	�T������,^��{f�U�%�|ov�IR��$�c*��h�A�����㮏	�nʝz�q~�6�������"ğ{�k���Ϻ�Vx��U��Y��Vg�MW�\��*��b�w4.��yqt�𬑺���Ȯ\G�L�,�em��:n�%���:�4/u���-����+0��
�G�g��~p��$��<��+�&g��^��:�]m��P
F��?l��	�������ţ���_���n:v�u9�s��7]��]`člM�=�]��ޱ�]�dk��߶�a����:��E~�'z�\m�B�+E�X�\&��w���Kd���IS)�F:�d����w�{4�)�����y�u
��T'D��v�:b�K���nX3���{��Wj�ut%)��_�����B��:6�I˘�����,:Ɇ¡���R�(ч_M�4���Q��j��n<��v4t�d�]�������yf���8K>a �_d�O~���@>��?�u���BQ�����ηY�ux?��t,'�+��	��&��PU��i�U�RU
<��K��3(��ZC�'�EB����.\��@�Nk$";�Ȱ��H��E\��G%2c$�T����O�u6��׃I1�5�]d�}凓���ZW�k]	�7�J�"�!ߘK6�1M����_��I�!_I���\韺��Ā�����邆�yA���
[ �ˢ­�YF!��|�t�a�J�ð9aa���7���Q=<��A[t!D�������~�!d7�qDpG)�<DM��۔�E�_��/Ǚ#m~Z��};�K�؆v?"/d�Q�s�����Ro54;��u��VJ��M�WS{�r�~���~���.� ��o���҇M$��13?��}�@u�n>`��������Am�yO!w\�->a� 'V5���o��m�׳%KG.��T���{�:W~���U�<OM��`o��|B!�?�$�jm�:[�Ԙ�e�n�Z�������}��/�����i�Π&�-���E��f(���4IG�(�Ǝ����� �����:�&{,���h��a���[��F�1��L�|�{{_��0;�ǜl/|rBc��i
9v���Ci�w0����sj��@XU�_�kn�������,L���rY�"0�d���ܮ
�W��u������d���oIH^"���������R�ބ��0��V�XRG�{bB�-�d5�"DO�+XlxVHYEB    fa00    1340NB��S�9���F\�a�?�zꪰA��
�M�Q%�s1��Q	0��@�1�W.�8�D���c��Cv^Ҿ�P�XOaM�!Hч!:X����H���7��p�*�Wڈ��}��\��8� ھ��s6[�P�wp�>u��j:��=P�4�j�������9H�=&{�gzg��nϔ"��}uxZ��rue���=Q��h7M�e�<f�sէ�hh��mY�ɩ.6�W�?�z^m������3y���(3��OC��1.���ﾯ�;.K ����t]���X���Q)f��Y��N�T�#�Ģ���&%l�*O��YUUV�-�y�g���P�pʊ��%I����zN.!��hz$7	�)��n����y�����0Bߴ�͎v&o<������ek|G���~3X�-O�"^;-z������Ȍ��z��W��:&�t�s~z�M[�Q�h�^���@2/���3(
���&�)g�|L���dg���Z.oC���L��aSWl3� �3o*��l�O�a�:�~5�A�{A1p�b���ة������ی	����7-q�[[`.�/<�B����x�F38~��C�n��V?�zͣ(/[�(��'Q=85�|d���H8�2b��D@/�Ĭk����#�:���#���i�N�B�����孼B���,N!.�P&$L��=�9�}g���\��VĄ��"PUBF��5 �N&DJ�^�r�lA�����������ߧħ:&�	:9#����.�:��)�U~)5K�#���ˡ��w0���K�ab5����7��O�k���`i�/B��3^=j>�«�e�EM�N<�ݸqA�e��'��g����rt����i?e_���� dl՟����0���c^�H�����ME&bf��̝��Eb^����W|[D&�����f�)�Uz�0X��h�u��s^�N����7
I(�,
�r'T^7Y��k�Q����,���ǭ�'���!�'x�z��G��qN2z4˥��<��w&0��`"�dp�n��z�$,%��M��������1�����G�i<B(n�n�{Y�g�;�\l!{�s"���F����x�(_�l�﵄�-:M9Ul��P��D1�)���o����˟����Z�r��j��]��z����+�F�������e�-���ڴ�5yΨ,��o[QZJd��dL���
� J{6k�
?��wʮ���R�B�_���r�"��.��8����q����a�;7���#L*v�u�d��m>p�W���)��{#E��7��J
�8E+�sO�W7��u��W��TN��a�&�f�f�|f�$�)t� �������%��b�mq��c���N�I����%��$�ُ�X�ש�/<��m�� �'�x|�5<�2���"���Ό�����!%��D��Y��.��+�1Pm���6����1L�2_�i	<�  v�`�ə"�&���k��+@�h�6�;��H�(�Z�;a��0K��M���f���V��:<@MBC���v瓃��� yG���;H���OZ���~�`G����d^�}.���w�p�Xz�A�&����eʀ��@�o�l�G�?�ѣ�p4����u�f�\j��ƦM@[#1��O�nY����H�x��VhR�њ���{�}��.f E۰��PƬn[8@�L��reT��w�Ĵ0;��	Ӱ4���i�a����v�K�C\���bg�Z�xT�f%�>"�#^Լ��[�~�	�ev�(�_h{�t@+:$e&��Vb,��u5���H��q���R��~%�Ι��.ʥ+�Ƚ�PbW�>���R+Y_x� V�����2�w��H�/ޭߕ��x�w�bf��*]YH��w�M�7l�ŉ~[ݯZ��g�63���9:Sa��g[E��_^�-�f�J����#b��59e>��&6y�T
����{���˚?�vd�?P5��?���w���⯼#�� �u�G���@�)�O����	d�w� �JgD��&�Ή�8���N�`�{��^�+�;��d��y�D�����ֈ׬?�@�̫�I��?!�ǻ�yA"����}�8�U�d��DFrE�5p{�ճqǻ��kj°2b����/E��$V�����r���c�L�]`< �q!�����4��8*�an"b����&Ou���=���Ka�B����0���]��R�Q\�8�R���\���-$X��7H�D@�61�C����b{w"E�f���IC����x�?�G:JlD��Zt�M�ӂ��;a����rf��M6v��!�9�v𬁨��ph�k23��	T�������B�غݯ�d%��ǎ���!&\��*�*H�{1t�N%��Q�vFqp��Б�8���}���J=_��Ҝ�]Bo�3#���;��A�7&rO��[��'{|��Cዊ��|�ɼex3�"JkaQB�]�UT�^p}W�L/�&|��.P��6+yl����]!@;�{j�\��
DnS��D��G7���.'���Ѱ�D(V9o�ʱ�c���gN� ��Z���O���5p�S���?�'�k5]qfNa��нL[��4����I2,4�fi_'}�����P�/A9id�d.FK�\m�N ��س�l�F(0��}*O�]`���컊^���d�f���+�F��+�'�}EO�1���x��A��}����r2l��Q��,��\8~ו�n��~�k���w�ܣ/���״-��D~�<��w|>,P�]��⧻%�Eќ��ȭM���*4 ޺�U�ʏB�q7P��$��w��P�x�ݟ44��Q(4M-��M��O�d���;�X�w��UF�^�]���T,�Qͧk-�U�ڃ�w�f���A!��u��zlA$`<��n��P6�
�q�AB
�?�������_�4�ִ~��$Pn
�5+��Nr�'g�T_0��z�vӗ+n~���G�����Q��VD-\�/��,v�@KN�Lk��c����͡o�������n�1�z~6U6oY�B=sbe	+�V����ț�^� �vG����ZL&|�������oҵ֣� ����jUP�@��q����]��lq�Ҝy�z��[i��B7�=s�(Mh�]�~�$�-��ø�]��̸�������U� zUb�h���eo�g�V`��݋gC�o�6�)gܒ2����E���)�h-�)o��D�A-��!����|�@�>o�&�U<���!�ڂe�Ǆ�L��c�q�k�Tj�T��)O��?s��ɕzb�c��x��o�G��/ۏ*?�+~1dKY�)Ι�Ƥ�>*��lJ�z*{���v�= 2�+�2�y���N�:dk�[����"�qY�Oұ/�!��2R~�tI���bD����v0��x$s�u�.	QS�x���U�_W��C,�2Q��� G��-_:�� �<�^��?$j�`�(I:�'�ũ>���ZL\<��IBFb��u+'2�i�#��q��/�Y� ��8��EvRV����[�2��KO0ŀ���H>$��}~�h<����W ��6�%����s�����l:�ٚ�������V+Q~2X��ʩ�6������G�-50�p����Np_[�0%v���0#�Su:��: TU~�z[�mѝ�L������L<Y�!$�%�g}�r)"�B#�Zx����=�c9�λ�&\ke��ˬ!�!Oz���.�����9q����N�k��e�%�A���1S�vI��������2����[һd>��c��V��­5���(�'������&'>A[Jۖ3��b#|T;���oǦz}��%@�����ŉ�Ig�d]ue���e���?v<�J*�a]y��6�*݅��z�/}�9���&��d��>�b�x�K������o�/fp�o�©H��J��+m*��!�hd��>~��2��e���P�	�v�&�^���:a�nB��V�8^��N��r�%O����}�����	����6��+1>����'���CƇbO�$$N�Q��?�{�����0�q�v��V$�f#�4�P�z�D3�|aň�̜��\��&�k��'�˞SX0���Ǜ�3���O�c�$DW@W� �F?�N�;�'���&��Q��v׺��CTf-�➙��,�>���l���O�ќb.D,��ueE��ԯՊ{�s�{
��7|�hۍ����ɹ8`�����q�-`�[��v�k�h�.���9�ءB��{ �^EW:=E��;�M�>�7�F��cM�7Y�9z�Kk����_w������)�gzN��I׼:��R
�mB��D�՗CiY$�W90�d�QQ,�a�ny{��4�[}��@[�i8�Лw#���3g���OHH�@���Y	�?z��F=ґ�RK�M?VI���ۂ���̶x�s�/�'�1�%�*��|}�8=�8#�PQ�\W�g] ��y�p�%��v�g�����!T����0�61s��C7׎��d�����@6%�UyV ����KN�M܋#Xb��j:�x!b��_����\�;�\�Tt&��=UGŐ�S���������C�2�ҽ.�&vu3�w��$tK��*v����\K���Ϟw�U�����^U>���ץծ��t&]����w�����+�yŮI&�&�cj��KLb����IBm��nW��\���>��d�&��eH\v-�����]�Q	:x? �)��I�ѫ�Հ�i-�+�eb�c�z��6����?��@U�הz(�o�z���UH�X�׌�&y�bi��?L�L^�ql*:����g�d\I`i�e�+]]!b_-�b�ɬU3XlxVHYEB      e7      a0�Ԋ�����&��bJ�42�Zˮ��"���,�1��ɏ�8��@�vO{	��K�ky`	Q��z?�>��5�G����1�����k��jj[g���~i�@��x���Y��|Ŏ�H�2&աj����T��ۣ�[�ԟI������{@řs�