XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���!a`���H@�e���=�S݇���t�C��5i@�J��
��۪H��i�\3��Gj2�{ͫ%�pt��N_����c=��j����ZO k�3��8�LSs��k�5�xa�{"�5Y�����kv�B�����GI=�����,?d��o��cn��ܻ5��(��pۺ�Y�UZmzDCK� ,��7�j�%o�c-OT����������D�/�@Z��Z<R�\�O��삐�b���RU.��[\���X�6%Tt�ĺup\�k���´�E@����i��+�ǻ���'Ux��)5��:��,��_�_U"�Q���eI�$|NW��E�눝=��?�}�g����0���E.���G����]��ō�W	�}�9 �_J��)��£�Yۤ����^�5�*��Ed�����5�C�2(
�Ȣ(t����e��b��fև2�M��1VS�t�E��[�0Т�;�#Ô��B7��R�&�޺b �<6Z�f�88;�"I��.kuA�;����az���-�O�SZ��"�xh��uT<?�ny���a�h;ۣ��ZvTN�M��9�(k:+���V��J����/,b�ŉ�����ؠ@
��W�/4e��v�:7�
�� O�!�n��DnX#�M+��vX�8H�pʄ1_�\^���	!�q�Zm�g! >z��� ��H`�.��LqoV����{
=��(6�ו1��^h�#�wA��-���OKK,7���-��V�L��/L����X5[m��XlxVHYEB    fa00    1950�D'E��}��/
λǷ���5����=���E.���s)"TSxD�GxY���̘��d~�;�k<���3�S����ȣm�u�56ʂ�OL���?'*rˏ�ü�oɯG�Xc�U����m��ē�����4���̷2:pt�5e�Do:�C;U���(G,���?Go��b�ꕐ��)�Mϻ��G��o���ހ�jOV����4����� J��;�W->A� �"�W�����^��X��I�h�+�)󇳜t,���jZ���k�ږv�1��?�e�,t�Q$�(������	��x�ZƟ!����&RR)1#*S/��I��nPs� �/�.��1p��e4���j��\�C[��6~�8<��4���[�qUͳ���t5�x����o�7��pP��7���8K\+ZԍT�Ϗ�u�jp���A�[��8�{%cb��yΩ`�Dj4f
�d�����!���:Hw������X�9D9��E���m	���Hp���*rQ �3�mo�d����+��~����0���������َ�޽V��P�wʾ�l��!�2�%���sy�T)-��������`���V�(f��D��.�Jf%ٍ�� ��a��Z	T�� �Y�墮�
�e߶�j�h:�ֺf�� >-]�i��4��e���� ��4c�k&�w]�5����d-�}�������-� 3򦼃|T�-r�#�����G�|A">8Pu�١�z�&���Y�����}�l!*�}6���������_끠����hP	҃�<(�[�얤�h��g�q�o-�Ni�nE���g�3l\�8�k�w�C����_g����
�t<<Mr�ϐ�zC�;�����W����F^��ơ"�~�_�za��4��N����u���?��0�|.�L�m�So:h��o�ƼaH沝�W��bh��w���4)w�"##=��+ȏ����.L2j���ϰ!��o�]8��r���G{��z��?h��^!����~�:k�49������w�Ĵ��kZ�{��Y�*\7p��Z�i����\T2׬mX����?/���.�}�&F�ےȧ�pnNG��z�a�y�J�[&�=@Q&�8(������X,�puXɚ�+w���p�Kkf2㑦w��;&�/K٧��=*^�^1���OH�A?1vI�xwf��1P���T��A�C2Ւ�z��' �C�Z�HR0~��B�&����QJ]+�DS��s�^!q�ұa�{=I'K��А ���jmҕ�Kc�^�I��S"M�FFNO4�F��a�I�#��u�iE�����B��0�`G��$�4���v��;,=�w/v�k疀l������E��c�-9�B�%��R�l0uh(dg�<���{a���X�ų˚�������q'9��>���,Q���c5�� R�}����hH���	�.w��X�򎛥��R��&(�@�&G!f1� �L;�s��������ei9����������`����4�� �g�R�]��P�?��+/�{�O�"?�[DPdҋ���Ӟ�����@����Z`���u�B����*��@��t�+t��!p��=�˿��msb� 7�w;=�s0e3[M~ɰ
�E�:��7	�# -� ��}b<���V=�"������|�1��X|��M�7�aq�P"�Zǘ��r�p�O�W/Ou�/<9�òB��ޡ
G<�Sn�� ��[|!q	�-QG�l�������O"�B8���7��٣C|u���v���DQ������� "4��k�����7�YJRż���G���4�Bo��_b��q:�G@���� K	�^Aɼ�C�V*��,��31���c/N �������x�hX��zZ�����ë�Ey��?(��i ���:�_�P��<&`��b��v�����ʟl�&S����Y�Ir|Q�臽s6��s't��1z�OJ�8�i��>���i��H�3�`�.d���,���\T+���дV��a_�7�v����YX�#�0����)�򻻇a���~az�8��v��:�
�O*J ĕ�S����C?��R[%!�m��<�w�5a���$�~��`w�0��0���^m���p�X�S��E��n��HL M�X;u`����������j�G%C�Ԟx�Df�L��9�����2�����)��,��='Y/��e�*h��I"(����o��0Ѹ�����-݌_��U\��,���4�UݟG��.��b�)���p�E]�f��R�8�������]�8�z��z��P6tt�\�(�T�p@���K�@O�U;Y9���ye��6���C�>R���#��#�~��]����Uv�������K�5
���we�^4������4ٷU����#G[{ex(Z9�Ya9���dl�[5c�0��4�b�
?�:���S���� �E	������������>e�v)[%�/%�ee	�ћ�h��|'�uUp��$!��Ds���{u���t��#X85�"��+������N�t��e5Ӫϭ|���0�v��oB�$Mg��K�o>F�o���7!���J�Jj "J��Bk{�yM{��#]�4���_+�ގ&R�h���x8^ig��IO{�@�����d(�K`1�����ߕ����xj��A"�۔`�k|��X����n0��鸢�0�vB|�W��i�z$���t7�[��i����pz��Yg"��߉��DǪ����O��0��pIÐ�^�u�0�\�淛�5�YƅAp���vݏ�)l�f��bJ^�T6<���/� �S�ov�& 5�/�Lv�W�'�u�=�)��]RN�C�q�g�o�$��S'/�����G�3�eNz�� ��>`>2�)���8���l̖v�.�h����D�z?ބ,���oQ��-]������[��D��/,i\.���G�G;FNa�)���[IWK�D1?�N>�����9B)y.����A�
�l��/aW�d��!������RH/T�H�`Zw�H<��~HzѾTKN��c/q��[�y�[��Y�d����+�+�%��&Ku:�H����^�S���,��O<1��A���2���>*�c�;���6*���_d�l��Ћ�V����Vm�ޙ_cރ��۟�4g}7M=��=��.V��Q�Q���؏�]9`�*Y|j|	���qJ s���dQ���&#�*@G�fmu�\so�df���BqV-�.��_����鎋*ש3�X6:g�x�haXZ���.S}��:hG�z�����0L')ߑ1�(.y����}6Yh���]�8�W[S<�(*!]�/!���/ӈ˖�tBQY�Pp�kL�8�~����|��|��޿9�&�go���>��$1Mo웍W�ڎ��L$l��V^T�hӃ�>;5�5�9�̹�?�zgah&i	�Rc���U�K
�����~��7���Y}���^4�W8b��m�:�����}��e7�vua6Ǣ�>��?�=��z�`M�����U�: v*�@��'��#OGq )�%�2C 
Ok:m��s+B*�;��U[r��p��9G�=_���l@c����@���;�\A�o���Ʃ����Of���a)�&�����?��Ô���$o��ǹL��.����k_v^jwP�s#���LWIEf�t��p.}:�+� �2lE�˘C���;R�͘�H�|u:Y�R,�Tz���5JvF��� o�g��~"p�E�������� `RZA�r:�ub�54u<� ��:���B.��1�vZ�]��y�gUEGZCI�-�� $��2N�٣�s�IǧǂV/ęӔ4h��-�
�:جPK9-ܦY(�毆���G�p;���O��ʞ� ��ߥ'x��U��wꂌj�֎S����|u'�5U�������L���f�\�
(FE���o[��c���~�hV4e�
t)&w����m�\����23Bwoѯ4��	�������G<��ҳ�OU헠����*����r�������pujN`p�Xj��\$�|�1�	)���73G�P>i�"�2��R�R�E7)m��}�˄���pV?Z	��F���4�V�G6^+B[�����Jʬ�13�E����`�HЁ+S5�3+�uXm8�8~�{Đ=J��q�(zS!�VJ���R�����RdyrF��+�IT|���]� ��J"���1?�Wm�����2���)�QTw��_t�\��fNw�g��.�ܾ�@�Z0�ʝ�o�&�u�E�4s����֊E+0���N.rsZ�$�z�p����OW¨��`?�uIz*����d����EHk�H;u{���"�����@�a�-�ڻR��_ϧ�B�w�a����0�;R�� G���RhE�GW��
*�9+l�5��Ɲ?8�:�	�&+��"W�m�z�jw݃�
q��%�4/{wx�1@�pc��3��m>G�gxV�������vc� ��s�_�Kk��M�y��NkX:C��jH�㭝u-�)�݅+8�Ѵވ$� ����u��TP��Gz�\�vX7��?��t�^8�<��f��#�G�j���wA4Slx_��J�jk���	�+�)��\No[���A�m9~-�<uZdx�--�R���jN@��<���
L�Mn�j?��d�ey�9J
�~`^uzׄ���jK�5���[�zWi��ڃD���o�Ԏ��a��?�&�>���D*�%��{��b7Ձ�/t�lUr�H�1@�C@am��ś�%
I�z�/�B�8��]$��T�q-0��j��ﺀ�3�}�z�e���2gd��H~�����\\Di&Ǖr]�C6.M��S뚺�~|����|~�و-8䟑��R�A�4y�T�����<�edY�j��VP�f$�2��n��t�f�z2�Tۜ�������~K�݉̿HO���G*F*��A��W Ao�~�vti:�G�&�Vi��q����K:+��\r����!~,�X�Y��T�����x�q�ª臨�@$��" O9�g� �L�-3��3��f%L�D ����f(D����+s���!�JIG�H>~{$��i�u���U�1��Y6�_nn)uD������MA�z�)��|F}���z��V��'�����@td��u`.sԥeȈ���	~8��?�I|p�]�_C=��Fƃq]�3�}�@-JY�(�H7�ݾ0WL'��#G��K�TbD��Fh~�r	���"���M�i���/k�u@'f�5^�U�Y�o�,1�(:}iX�m��a�����X��j�C��2��ځ�=r��\a=�Ā�e�$��^_܉xsA
�"(� 
 4\����x�#�%�A(�����v��|R�h�g�Ǳ���qe	v��ߨ5[��4��1&uu������0A �nn�'/�\Ð�B{�O�T�h�^2�~[*)�K������H=k!������ ������[�}	aa���`("�:0����D���a`����S$\��²�c���v�G��\��"�zUDؑ�h���.�<`���0�:ÀS"���=e�Kx���t:����P�r�]Ǽ���ۓ����+���?%�ƒ!o4�g�@]��XT�����3x<� ��ek��XI��
�8b&��KI�.��}B�%`ϫf)p���ެf���ё�7�k�RW�>߃%��b��"߰�Q<���NE7�`_�'BБ����p{�f���}5��+��b�*"9����[�(�0c�"�;(�f��A!�x.�sR�Ք԰V�.3Αnk��n�����{��q�Sb�w��#!��$݈; �h���1^��o��q��+kU�W��T�y�E�qD�2D1Ȕ�U���H�CA���6-T�,�υT^����&t��l���t,c�K	����G���I|�T߇E����UD�A`�r�U��@�mȧعY�Fw��)kP3����P_E��wQ	aI��x7�?6H,�G`�-�eʕ����I�!P�N/%�����yFdTl$�֤_ ��P����S�����3o���J�7���6�	�=�'�]f0M[ą[(��rˮ:@#��b�ǻ�2�Y�4�֤dR�q��/rh�.����h��y�-!+��]��Y�D�`i�����c��g��-���G��Ħ��� �7�`ȥ�W�D�\>+B�b��އ�IJm2��n�o%30�/?��GѶr_gY�sUR�qk�|爿��)Q}�{�öq�R �	$g�!��u��#c�Q��t\�1݃�d�T�!2B��)��h���t��A�&B�!@�����zf�t��۲o�%L��"�/?��U-�ǆ2��޽�������Y�5N�ެC����)QvrA�@�%ěXlxVHYEB    fa00     700�e��2����~ňDe�ʁ����D�H����\�rC�s˲�)+����8nq�Ku���с	k�!�V����v̚nb��f�<Z�vG�g�O-�a�7d���R"֘jY���ݔM-�>�����B<>����y��VEOr�� �W|@\ua�C#�c�\��rXo�ȃ}��48@����sl�;���8�zO�%sv��ұ���Jy���M_�!�^�N/�jՃ�yI]���[
�+�"�oCH�V6����P��,!y-�M�q�gH�l7L_/t`�I�3�ɵ �X6���,n�� �C?at�"C�T��4^t({T�z�A�L�9z��i"�j�0k���y�b���oMb���^ɑK�샏�1,�Rnq������L�f?�e�;�o����u�C�����|bT}�}c�p�iS���n��*����m��)��^�c����x�l]8��&�d���̝4l���[r�z/І�k�P�����x[�ASI|^����*�z�5���"&�9,~��YM�.|*�^�	��|�G{��2�/zW�^�t���;�o��`�$����;$XN��̜�~P@��n�/��
"�r�����?޹9~�s���������i�.���xbץ���\��o�$! ����}l�3#�D���C�
�j��� ���ԛ�>�. ��|�q�0;�*��4�Yx	�����$S�@0����b��DA x�rw7&`ؐ$����yF>�<�T��}��T�Om��S.c�4nL�aG��^DZ��'R_s���>����h����3��]h5^�c(��D�X�=m�����.+8�7%%��^���Aa�S�@��Y�^)!�?ӭZb�qu��z���� ��E�_?F�c�?{��J[^e_����e�KsM���%��N௼Yưp�<,l��
Sc�5ڋ�,L�'�|i=���̪Kt"j;����o<�Q�U�Nw��hQ�t-}�i�5'���h�%��?��iR�@�2�cC�Dr����p�m�:{�r}��"TA�ʂE��j���΍��w�V`��8�{��4�(ߢ��h��g���]5��`��d��9d�ėqǸ&�(�y��\���x"i��{�������ݏ�� ��9���f�G,.��ᮟr�"1�h�F%�E�>�Y~�W�H�W�������CiF00}�顏Xk�V�nX�LN��'y�5��&磲[DsG�>��R.CMe��Z�����aAC ��P�ꊼ��U~��u֏��O�e';����$V
�1	?n�b�Sb'�+vO��,�Ʉ袏�98���-q�B�]$ƕ�g]�ѭmڶ�Ɋ/'��E�]�͸˄{�ȶS�`|t�����	��s�|�l�!5����H>=�{�lz��:b�^�%�c��YZ`�*)r�0�O,L�_��`�8$���b�Fȹ+�`թ&�Uޞ��_t�>|s҃�dc[ �`��	��H�ފ���i��+�Y�UOw�sD�Z+�ؗ�?�� ��H�,��ڬs����m~H�.ZQe���M*EL�?i�fa�2�WDeQ�p�=I
�睇�.JCc���:�>�O�3�2�J2���ɞ6(�㊄GxQ)��hDř�-)����qb9HM$������5YV1���!8�a�i`�r?[�y���,�eEo
)H@b�*�'|��:`Cj.T|��\tD&D��(�_�--v����"�~S�lB��0N+�� ,�Q���o�*�I4͛x>>�͝a��N� �����j���'XlxVHYEB    77da     a60�� b�q7,��6X��Fs��jOn��y+�b$�g����*A�sxaN�P��]�������UH�X	n���=��<���0�p)�����bJ��M^����2ƣ-yھ��c\����Gh�c*s-�~}����fN�Z�d��~�!��s�?#e��OM��q��Ɛ
�ѫ��@�S���1fA1^~|�C�h����r�����;j��x�QyuK f��C�����兩|̌^��f�B	�(
��Ǧt1܂.!���33
/1��h��y	�N��7ϵu��Gn/'��{�0��<�2°��D���\��1t:OwBw���uy*rX�LÌ�"��J%#9�����衠Ǳ'����Н��M-���BH!4HM��mq��A����=���)w9��1�w�{��|�n8���7� C�7,
�[�x�|z��ֵt�1�H�}m�6B?Л�[A�A�0m��X�L^��2����G�2������0b�Q
3��n����/�Y���5`����}\}�$���+ƶ߉�� br7�3ɺ�jf"f��Kς��i�۵�+I���úF��1��E��?
��4P �+��;r壳E��g��v��:�EB�A9�����)'�Q��S	l)�D��ń�U�-h��D�G��F�ȩ�;��L	W"�Jo4J�ou��U�o�I�8˓! �W���/�3Lg�:M�uk�DI��Ahl3x���ת1�4ۚ8!�۲V����e���UuS$�ˢf@�ιT{��]�K,4��lˀ�V�a�cQv�URς�H�t9�v���ˑ����+f��̂@B�n[�Q2��"��+K)v���k67Xk��^���'��������~�����:P��F��H���t�z�C�T�k8���ُ���޳ʝ�6�i|��6anB�����̐�h��+Y[z0o�8�.h� �[���VY�r�+:���5���r�/U%۝;����g�95J� ��R��3��[5~�T��%@F[�X�8��='�� 9f��i�LH�CXU�??�3i����dS����	��cL��4_���B-�/�чWm�v�	�1_��/�dV���l�@X���� }V����)�}���D��;���,s�&�6W�⪭B�b�� ܅��?^^�|a�3w�d�_}�8,\q������A��=L9�/�AKs�ꈰ��<���g��_�Xl�ߦ� n��%�l�[s��l�/Ux�?�7�7�R��d��W)��e@�62����U���b�:#H�vy��R8\�Ʋ�rf3�S�f��ܪ�%��֖��a�
���Io{��'X�5�T���h9#1I����ԉ���$nae�.�/�~4=�m�e���X�5����>�ԀeVg��."���R�Z�L���A<����5 `���%o�l�кx�d��%��,C��Q�Ʀ���倃�b�5���$�!�{;_��\��՛%sFc�4xA�\�O݃�Y�d���FOoW͜م\�U����~�	7��\�S f�:�W2��6�Z86���p��`�D��eh�u���b�48Dah�y��9�-̜�~��}�l��{rD>����F��W�����]���ځ�������)�D�,j���e7�7�?}��{{�&^���%��T���j*��g�t�$����K��6��%^�w�a����%��]�6c�%s��0���i�<�w��A%`���� $���;����: ���܈��
��ֱb�i�q��;������F���ӔLx��k���yt\��M����d�Qx�����/�ޠ�v�Þ&7
۟IjG�����ddD��C��-��XUCd�����(�U;��|W ʲL��=�-~�$!��S�<���^҃<�n#�O�L�=�ɦ�n��?���i���S'E������j:$��ѯ�;E�*ʤ7x0�8�/�XW_M��h� �A2�ΒH���ß���V!�ӱw0�nd�v�8A��� >�PkXm��\�A��ӯ�ajQ�B�$ji.rW���&�͕�`_-�t�.p����< ��>({q���'�_�̠� ���R`��o��dd��+)�!��y!�U��h������nr�dZ�K#��?�Τ%���"`�������^��\_ߋ�XxDP`�P�LT[��� Dx�)鼧�-h*���	� ���A�W&i���z�.��	�
�Ł|g�hb<�V�+���FQ=���UTs���8��s�Y�U/��э/�8��e�*��`�-�=I����xlSe+����\�
ޓ���=͢@��X1>�w�a�8n<�tKrg��G9����*,�X�t���C*�y%P9�H���y�F���O����=�j�`�],� 3pㆄh����@��&Xd�П��flh�$�8 ty�ǜ`1取��6���U����?$�LC�z�bu=����6�Y�4��%3�6�0@�8���|@�Bg�� ��w��A�+��� �&}J���'���yl�AR��8�{���:�����d.b�N��&cR8t`�����F'���m���nm�f��^����x���=�3zյ T&'��'�K���Fj�恾�U���gxA�7Zsw  �"